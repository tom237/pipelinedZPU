`timescale 1ns / 1ps

module memory(
    input wire clk,
    input wire[3:0] wea,
    input wire[31:0] dina,
    input wire ena,
    output reg[31:0] douta,
    input wire[31:0] addra,

    output reg[31:0] doutb,
    input wire[3:0] web,
    input wire[31:0] dinb,
    input wire enb,
    input wire[31:0] addrb
);


    reg[31:0] RAM[8192:0];

    initial begin
        RAM[1] = 32'h82700b0b,
        RAM[2] = 32'h80ceb40c,
        RAM[3] = 32'h3a0b0b80,
        RAM[4] = 32'hc6c20400,
        RAM[5] = 32'h00000000,
        RAM[6] = 32'h00000000,
        RAM[7] = 32'h00000000,
        RAM[8] = 32'h00000000,
        RAM[9] = 32'h90089408,
        RAM[10] = 32'h980881a0,
        RAM[11] = 32'h900a080b,
        RAM[12] = 32'h0b80cec0,
        RAM[13] = 32'h05082d98,
        RAM[14] = 32'h0c940c90,
        RAM[15] = 32'h0c030400,
        RAM[16] = 32'h00000000,
        RAM[17] = 32'h71fd0608,
        RAM[18] = 32'h72830609,
        RAM[19] = 32'h81058205,
        RAM[20] = 32'h832b2a83,
        RAM[21] = 32'hffff0652,
        RAM[22] = 32'h04000000,
        RAM[23] = 32'h00000000,
        RAM[24] = 32'h00000000,
        RAM[25] = 32'h71fd0608,
        RAM[26] = 32'h83ffff73,
        RAM[27] = 32'h83060981,
        RAM[28] = 32'h05820583,
        RAM[29] = 32'h2b2b0906,
        RAM[30] = 32'h7383ffff,
        RAM[31] = 32'h0b0b0b0b,
        RAM[32] = 32'h83a70400,
        RAM[33] = 32'h72098105,
        RAM[34] = 32'h72057373,
        RAM[35] = 32'h09060906,
        RAM[36] = 32'h73097306,
        RAM[37] = 32'h070a8106,
        RAM[38] = 32'h53510400,
        RAM[39] = 32'h00000000,
        RAM[40] = 32'h00000000,
        RAM[41] = 32'h72722473,
        RAM[42] = 32'h732e0753,
        RAM[43] = 32'h51040000,
        RAM[44] = 32'h00000000,
        RAM[45] = 32'h00000000,
        RAM[46] = 32'h00000000,
        RAM[47] = 32'h00000000,
        RAM[48] = 32'h00000000,
        RAM[49] = 32'h71737109,
        RAM[50] = 32'h71068106,
        RAM[51] = 32'h30720a10,
        RAM[52] = 32'h0a720a10,
        RAM[53] = 32'h0a31050a,
        RAM[54] = 32'h81065151,
        RAM[55] = 32'h53510400,
        RAM[56] = 32'h00000000,
        RAM[57] = 32'h72722673,
        RAM[58] = 32'h732e0753,
        RAM[59] = 32'h51040000,
        RAM[60] = 32'h00000000,
        RAM[61] = 32'h00000000,
        RAM[62] = 32'h00000000,
        RAM[63] = 32'h00000000,
        RAM[64] = 32'h00000000,
        RAM[65] = 32'h00000000,
        RAM[66] = 32'h00000000,
        RAM[67] = 32'h00000000,
        RAM[68] = 32'h00000000,
        RAM[69] = 32'h00000000,
        RAM[70] = 32'h00000000,
        RAM[71] = 32'h00000000,
        RAM[72] = 32'h00000000,
        RAM[73] = 32'h0b0b0b88,
        RAM[74] = 32'hc4040000,
        RAM[75] = 32'h00000000,
        RAM[76] = 32'h00000000,
        RAM[77] = 32'h00000000,
        RAM[78] = 32'h00000000,
        RAM[79] = 32'h00000000,
        RAM[80] = 32'h00000000,
        RAM[81] = 32'h720a722b,
        RAM[82] = 32'h0a535104,
        RAM[83] = 32'h00000000,
        RAM[84] = 32'h00000000,
        RAM[85] = 32'h00000000,
        RAM[86] = 32'h00000000,
        RAM[87] = 32'h00000000,
        RAM[88] = 32'h00000000,
        RAM[89] = 32'h72729f06,
        RAM[90] = 32'h0981050b,
        RAM[91] = 32'h0b0b88a7,
        RAM[92] = 32'h05040000,
        RAM[93] = 32'h00000000,
        RAM[94] = 32'h00000000,
        RAM[95] = 32'h00000000,
        RAM[96] = 32'h00000000,
        RAM[97] = 32'h72722aff,
        RAM[98] = 32'h739f062a,
        RAM[99] = 32'h0974090a,
        RAM[100] = 32'h8106ff05,
        RAM[101] = 32'h06075351,
        RAM[102] = 32'h04000000,
        RAM[103] = 32'h00000000,
        RAM[104] = 32'h00000000,
        RAM[105] = 32'h71715351,
        RAM[106] = 32'h020d0406,
        RAM[107] = 32'h73830609,
        RAM[108] = 32'h81058205,
        RAM[109] = 32'h832b0b2b,
        RAM[110] = 32'h0772fc06,
        RAM[111] = 32'h0c515104,
        RAM[112] = 32'h00000000,
        RAM[113] = 32'h72098105,
        RAM[114] = 32'h72050970,
        RAM[115] = 32'h81050906,
        RAM[116] = 32'h0a810653,
        RAM[117] = 32'h51040000,
        RAM[118] = 32'h00000000,
        RAM[119] = 32'h00000000,
        RAM[120] = 32'h00000000,
        RAM[121] = 32'h72098105,
        RAM[122] = 32'h72050970,
        RAM[123] = 32'h81050906,
        RAM[124] = 32'h0a098106,
        RAM[125] = 32'h53510400,
        RAM[126] = 32'h00000000,
        RAM[127] = 32'h00000000,
        RAM[128] = 32'h00000000,
        RAM[129] = 32'h71098105,
        RAM[130] = 32'h52040000,
        RAM[131] = 32'h00000000,
        RAM[132] = 32'h00000000,
        RAM[133] = 32'h00000000,
        RAM[134] = 32'h00000000,
        RAM[135] = 32'h00000000,
        RAM[136] = 32'h00000000,
        RAM[137] = 32'h72720981,
        RAM[138] = 32'h05055351,
        RAM[139] = 32'h04000000,
        RAM[140] = 32'h00000000,
        RAM[141] = 32'h00000000,
        RAM[142] = 32'h00000000,
        RAM[143] = 32'h00000000,
        RAM[144] = 32'h00000000,
        RAM[145] = 32'h72097206,
        RAM[146] = 32'h73730906,
        RAM[147] = 32'h07535104,
        RAM[148] = 32'h00000000,
        RAM[149] = 32'h00000000,
        RAM[150] = 32'h00000000,
        RAM[151] = 32'h00000000,
        RAM[152] = 32'h00000000,
        RAM[153] = 32'h71fc0608,
        RAM[154] = 32'h72830609,
        RAM[155] = 32'h81058305,
        RAM[156] = 32'h1010102a,
        RAM[157] = 32'h81ff0652,
        RAM[158] = 32'h04000000,
        RAM[159] = 32'h00000000,
        RAM[160] = 32'h00000000,
        RAM[161] = 32'h71fc0608,
        RAM[162] = 32'h0b0b80cd,
        RAM[163] = 32'hf8738306,
        RAM[164] = 32'h10100508,
        RAM[165] = 32'h060b0b0b,
        RAM[166] = 32'h88aa0400,
        RAM[167] = 32'h00000000,
        RAM[168] = 32'h00000000,
        RAM[169] = 32'h0b0b0b88,
        RAM[170] = 32'hf8040000,
        RAM[171] = 32'h00000000,
        RAM[172] = 32'h00000000,
        RAM[173] = 32'h00000000,
        RAM[174] = 32'h00000000,
        RAM[175] = 32'h00000000,
        RAM[176] = 32'h00000000,
        RAM[177] = 32'h0b0b0b88,
        RAM[178] = 32'he0040000,
        RAM[179] = 32'h00000000,
        RAM[180] = 32'h00000000,
        RAM[181] = 32'h00000000,
        RAM[182] = 32'h00000000,
        RAM[183] = 32'h00000000,
        RAM[184] = 32'h00000000,
        RAM[185] = 32'h72097081,
        RAM[186] = 32'h0509060a,
        RAM[187] = 32'h8106ff05,
        RAM[188] = 32'h70547106,
        RAM[189] = 32'h73097274,
        RAM[190] = 32'h05ff0506,
        RAM[191] = 32'h07515151,
        RAM[192] = 32'h04000000,
        RAM[193] = 32'h72097081,
        RAM[194] = 32'h0509060a,
        RAM[195] = 32'h098106ff,
        RAM[196] = 32'h05705471,
        RAM[197] = 32'h06730972,
        RAM[198] = 32'h7405ff05,
        RAM[199] = 32'h06075151,
        RAM[200] = 32'h51040000,
        RAM[201] = 32'h05ff0504,
        RAM[202] = 32'h00000000,
        RAM[203] = 32'h00000000,
        RAM[204] = 32'h00000000,
        RAM[205] = 32'h00000000,
        RAM[206] = 32'h00000000,
        RAM[207] = 32'h00000000,
        RAM[208] = 32'h00000000,
        RAM[209] = 32'h810b0b0b,
        RAM[210] = 32'h80ceb00c,
        RAM[211] = 32'h51040000,
        RAM[212] = 32'h00000000,
        RAM[213] = 32'h00000000,
        RAM[214] = 32'h00000000,
        RAM[215] = 32'h00000000,
        RAM[216] = 32'h00000000,
        RAM[217] = 32'h71810552,
        RAM[218] = 32'h04000000,
        RAM[219] = 32'h00000000,
        RAM[220] = 32'h00000000,
        RAM[221] = 32'h00000000,
        RAM[222] = 32'h00000000,
        RAM[223] = 32'h00000000,
        RAM[224] = 32'h00000000,
        RAM[225] = 32'h00000000,
        RAM[226] = 32'h00000000,
        RAM[227] = 32'h00000000,
        RAM[228] = 32'h00000000,
        RAM[229] = 32'h00000000,
        RAM[230] = 32'h00000000,
        RAM[231] = 32'h00000000,
        RAM[232] = 32'h00000000,
        RAM[233] = 32'h02840572,
        RAM[234] = 32'h10100552,
        RAM[235] = 32'h04000000,
        RAM[236] = 32'h00000000,
        RAM[237] = 32'h00000000,
        RAM[238] = 32'h00000000,
        RAM[239] = 32'h00000000,
        RAM[240] = 32'h00000000,
        RAM[241] = 32'h00000000,
        RAM[242] = 32'h00000000,
        RAM[243] = 32'h00000000,
        RAM[244] = 32'h00000000,
        RAM[245] = 32'h00000000,
        RAM[246] = 32'h00000000,
        RAM[247] = 32'h00000000,
        RAM[248] = 32'h00000000,
        RAM[249] = 32'h717105ff,
        RAM[250] = 32'h05715351,
        RAM[251] = 32'h020d0400,
        RAM[252] = 32'h00000000,
        RAM[253] = 32'h00000000,
        RAM[254] = 32'h00000000,
        RAM[255] = 32'h00000000,
        RAM[256] = 32'h00000000,
        RAM[257] = 32'h82f53f80,
        RAM[258] = 32'hc5c43f04,
        RAM[259] = 32'h10101010,
        RAM[260] = 32'h10101010,
        RAM[261] = 32'h10101010,
        RAM[262] = 32'h10101010,
        RAM[263] = 32'h10101010,
        RAM[264] = 32'h10101010,
        RAM[265] = 32'h10101010,
        RAM[266] = 32'h10101053,
        RAM[267] = 32'h51047381,
        RAM[268] = 32'hff067383,
        RAM[269] = 32'h06098105,
        RAM[270] = 32'h83051010,
        RAM[271] = 32'h102b0772,
        RAM[272] = 32'hfc060c51,
        RAM[273] = 32'h51043c04,
        RAM[274] = 32'h72728072,
        RAM[275] = 32'h8106ff05,
        RAM[276] = 32'h09720605,
        RAM[277] = 32'h71105272,
        RAM[278] = 32'h0a100a53,
        RAM[279] = 32'h72ed3851,
        RAM[280] = 32'h51535104,
        RAM[281] = 32'h90089408,
        RAM[282] = 32'h98087575,
        RAM[283] = 32'h8df02d50,
        RAM[284] = 32'h50900856,
        RAM[285] = 32'h980c940c,
        RAM[286] = 32'h900c5104,
        RAM[287] = 32'h90089408,
        RAM[288] = 32'h98087575,
        RAM[289] = 32'h8cbe2d50,
        RAM[290] = 32'h50900856,
        RAM[291] = 32'h980c940c,
        RAM[292] = 32'h900c5104,
        RAM[293] = 32'hfe3d0d0b,
        RAM[294] = 32'h0b80df9c,
        RAM[295] = 32'h08538413,
        RAM[296] = 32'h0870882a,
        RAM[297] = 32'h70810651,
        RAM[298] = 32'h52527080,
        RAM[299] = 32'h2ef03871,
        RAM[300] = 32'h81ff0690,
        RAM[301] = 32'h0c843d0d,
        RAM[302] = 32'h04ff3d0d,
        RAM[303] = 32'h0b0b80df,
        RAM[304] = 32'h9c085271,
        RAM[305] = 32'h0870882a,
        RAM[306] = 32'h81327081,
        RAM[307] = 32'h06515151,
        RAM[308] = 32'h70f13873,
        RAM[309] = 32'h720c833d,
        RAM[310] = 32'h0d0480ce,
        RAM[311] = 32'hb008802e,
        RAM[312] = 32'ha43880ce,
        RAM[313] = 32'hb408822e,
        RAM[314] = 32'hbd388380,
        RAM[315] = 32'h800b0b0b,
        RAM[316] = 32'h80df9c0c,
        RAM[317] = 32'h82a0800b,
        RAM[318] = 32'h80dfa00c,
        RAM[319] = 32'h8290800b,
        RAM[320] = 32'h80dfa40c,
        RAM[321] = 32'h04f88080,
        RAM[322] = 32'h80a40b0b,
        RAM[323] = 32'h0b80df9c,
        RAM[324] = 32'h0cf88080,
        RAM[325] = 32'h82800b80,
        RAM[326] = 32'hdfa00cf8,
        RAM[327] = 32'h80808480,
        RAM[328] = 32'h0b80dfa4,
        RAM[329] = 32'h0c0480c0,
        RAM[330] = 32'ha8808c0b,
        RAM[331] = 32'h0b0b80df,
        RAM[332] = 32'h9c0c80c0,
        RAM[333] = 32'ha880940b,
        RAM[334] = 32'h80dfa00c,
        RAM[335] = 32'h80ce880b,
        RAM[336] = 32'h80dfa40c,
        RAM[337] = 32'h04ff3d0d,
        RAM[338] = 32'h80dfa833,
        RAM[339] = 32'h5170a738,
        RAM[340] = 32'h80cebc08,
        RAM[341] = 32'h70085252,
        RAM[342] = 32'h70802e94,
        RAM[343] = 32'h38841280,
        RAM[344] = 32'hcebc0c70,
        RAM[345] = 32'h2d80cebc,
        RAM[346] = 32'h08700852,
        RAM[347] = 32'h5270ee38,
        RAM[348] = 32'h810b80df,
        RAM[349] = 32'ha834833d,
        RAM[350] = 32'h0d040480,
        RAM[351] = 32'h3d0d0b0b,
        RAM[352] = 32'h80df9808,
        RAM[353] = 32'h802e8e38,
        RAM[354] = 32'h0b0b0b0b,
        RAM[355] = 32'h800b802e,
        RAM[356] = 32'h09810685,
        RAM[357] = 32'h38823d0d,
        RAM[358] = 32'h040b0b80,
        RAM[359] = 32'hdf98510b,
        RAM[360] = 32'h0b0bf4e0,
        RAM[361] = 32'h3f823d0d,
        RAM[362] = 32'h0404830b,
        RAM[363] = 32'h80c0a880,
        RAM[364] = 32'ha00cff39,
        RAM[365] = 32'h810b80c0,
        RAM[366] = 32'ha880b00c,
        RAM[367] = 32'h04803d0d,
        RAM[368] = 32'h80ce8c51,
        RAM[369] = 32'h86d33f81,
        RAM[370] = 32'h0b80c0a8,
        RAM[371] = 32'h80b00c82,
        RAM[372] = 32'h3d0d0480,
        RAM[373] = 32'h3d0d80c0,
        RAM[374] = 32'ha8808c08,
        RAM[375] = 32'h70882a81,
        RAM[376] = 32'h32708106,
        RAM[377] = 32'h51515170,
        RAM[378] = 32'hed3880c0,
        RAM[379] = 32'ha8809008,
        RAM[380] = 32'h7081ff06,
        RAM[381] = 32'h80c0a880,
        RAM[382] = 32'h8c0c5181,
        RAM[383] = 32'h0b80c0a8,
        RAM[384] = 32'h80a80c82,
        RAM[385] = 32'h3d0d0483,
        RAM[386] = 32'h0b80c0a8,
        RAM[387] = 32'h80a00cc0,
        RAM[388] = 32'h0a0b80c0,
        RAM[389] = 32'ha880b40c,
        RAM[390] = 32'h830b80c0,
        RAM[391] = 32'ha880b00c,
        RAM[392] = 32'h810b80c0,
        RAM[393] = 32'ha880ac0c,
        RAM[394] = 32'h810b80c0,
        RAM[395] = 32'ha880a40c,
        RAM[396] = 32'h810b80c0,
        RAM[397] = 32'ha8809c0c,
        RAM[398] = 32'h800b80c0,
        RAM[399] = 32'ha880a00c,
        RAM[400] = 32'hff399c08,
        RAM[401] = 32'h029c0cf9,
        RAM[402] = 32'h3d0d800b,
        RAM[403] = 32'h9c08fc05,
        RAM[404] = 32'h0c9c0888,
        RAM[405] = 32'h05088025,
        RAM[406] = 32'hab389c08,
        RAM[407] = 32'h88050830,
        RAM[408] = 32'h9c088805,
        RAM[409] = 32'h0c800b9c,
        RAM[410] = 32'h08f4050c,
        RAM[411] = 32'h9c08fc05,
        RAM[412] = 32'h08883881,
        RAM[413] = 32'h0b9c08f4,
        RAM[414] = 32'h050c9c08,
        RAM[415] = 32'hf405089c,
        RAM[416] = 32'h08fc050c,
        RAM[417] = 32'h9c088c05,
        RAM[418] = 32'h088025ab,
        RAM[419] = 32'h389c088c,
        RAM[420] = 32'h0508309c,
        RAM[421] = 32'h088c050c,
        RAM[422] = 32'h800b9c08,
        RAM[423] = 32'hf0050c9c,
        RAM[424] = 32'h08fc0508,
        RAM[425] = 32'h8838810b,
        RAM[426] = 32'h9c08f005,
        RAM[427] = 32'h0c9c08f0,
        RAM[428] = 32'h05089c08,
        RAM[429] = 32'hfc050c80,
        RAM[430] = 32'h539c088c,
        RAM[431] = 32'h0508529c,
        RAM[432] = 32'h08880508,
        RAM[433] = 32'h5181a73f,
        RAM[434] = 32'h9008709c,
        RAM[435] = 32'h08f8050c,
        RAM[436] = 32'h549c08fc,
        RAM[437] = 32'h0508802e,
        RAM[438] = 32'h8c389c08,
        RAM[439] = 32'hf8050830,
        RAM[440] = 32'h9c08f805,
        RAM[441] = 32'h0c9c08f8,
        RAM[442] = 32'h05087090,
        RAM[443] = 32'h0c54893d,
        RAM[444] = 32'h0d9c0c04,
        RAM[445] = 32'h9c08029c,
        RAM[446] = 32'h0cfb3d0d,
        RAM[447] = 32'h800b9c08,
        RAM[448] = 32'hfc050c9c,
        RAM[449] = 32'h08880508,
        RAM[450] = 32'h80259338,
        RAM[451] = 32'h9c088805,
        RAM[452] = 32'h08309c08,
        RAM[453] = 32'h88050c81,
        RAM[454] = 32'h0b9c08fc,
        RAM[455] = 32'h050c9c08,
        RAM[456] = 32'h8c050880,
        RAM[457] = 32'h258c389c,
        RAM[458] = 32'h088c0508,
        RAM[459] = 32'h309c088c,
        RAM[460] = 32'h050c8153,
        RAM[461] = 32'h9c088c05,
        RAM[462] = 32'h08529c08,
        RAM[463] = 32'h88050851,
        RAM[464] = 32'had3f9008,
        RAM[465] = 32'h709c08f8,
        RAM[466] = 32'h050c549c,
        RAM[467] = 32'h08fc0508,
        RAM[468] = 32'h802e8c38,
        RAM[469] = 32'h9c08f805,
        RAM[470] = 32'h08309c08,
        RAM[471] = 32'hf8050c9c,
        RAM[472] = 32'h08f80508,
        RAM[473] = 32'h70900c54,
        RAM[474] = 32'h873d0d9c,
        RAM[475] = 32'h0c049c08,
        RAM[476] = 32'h029c0cfd,
        RAM[477] = 32'h3d0d810b,
        RAM[478] = 32'h9c08fc05,
        RAM[479] = 32'h0c800b9c,
        RAM[480] = 32'h08f8050c,
        RAM[481] = 32'h9c088c05,
        RAM[482] = 32'h089c0888,
        RAM[483] = 32'h050827ac,
        RAM[484] = 32'h389c08fc,
        RAM[485] = 32'h0508802e,
        RAM[486] = 32'ha338800b,
        RAM[487] = 32'h9c088c05,
        RAM[488] = 32'h08249938,
        RAM[489] = 32'h9c088c05,
        RAM[490] = 32'h08109c08,
        RAM[491] = 32'h8c050c9c,
        RAM[492] = 32'h08fc0508,
        RAM[493] = 32'h109c08fc,
        RAM[494] = 32'h050cc939,
        RAM[495] = 32'h9c08fc05,
        RAM[496] = 32'h08802e80,
        RAM[497] = 32'hc9389c08,
        RAM[498] = 32'h8c05089c,
        RAM[499] = 32'h08880508,
        RAM[500] = 32'h26a1389c,
        RAM[501] = 32'h08880508,
        RAM[502] = 32'h9c088c05,
        RAM[503] = 32'h08319c08,
        RAM[504] = 32'h88050c9c,
        RAM[505] = 32'h08f80508,
        RAM[506] = 32'h9c08fc05,
        RAM[507] = 32'h08079c08,
        RAM[508] = 32'hf8050c9c,
        RAM[509] = 32'h08fc0508,
        RAM[510] = 32'h812a9c08,
        RAM[511] = 32'hfc050c9c,
        RAM[512] = 32'h088c0508,
        RAM[513] = 32'h812a9c08,
        RAM[514] = 32'h8c050cff,
        RAM[515] = 32'haf399c08,
        RAM[516] = 32'h90050880,
        RAM[517] = 32'h2e8f389c,
        RAM[518] = 32'h08880508,
        RAM[519] = 32'h709c08f4,
        RAM[520] = 32'h050c518d,
        RAM[521] = 32'h399c08f8,
        RAM[522] = 32'h0508709c,
        RAM[523] = 32'h08f4050c,
        RAM[524] = 32'h519c08f4,
        RAM[525] = 32'h0508900c,
        RAM[526] = 32'h853d0d9c,
        RAM[527] = 32'h0c04fc3d,
        RAM[528] = 32'h0d767079,
        RAM[529] = 32'h7b555555,
        RAM[530] = 32'h558f7227,
        RAM[531] = 32'h8c387275,
        RAM[532] = 32'h07830651,
        RAM[533] = 32'h70802ea7,
        RAM[534] = 32'h38ff1252,
        RAM[535] = 32'h71ff2e98,
        RAM[536] = 32'h38727081,
        RAM[537] = 32'h05543374,
        RAM[538] = 32'h70810556,
        RAM[539] = 32'h34ff1252,
        RAM[540] = 32'h71ff2e09,
        RAM[541] = 32'h8106ea38,
        RAM[542] = 32'h74900c86,
        RAM[543] = 32'h3d0d0474,
        RAM[544] = 32'h51727084,
        RAM[545] = 32'h05540871,
        RAM[546] = 32'h70840553,
        RAM[547] = 32'h0c727084,
        RAM[548] = 32'h05540871,
        RAM[549] = 32'h70840553,
        RAM[550] = 32'h0c727084,
        RAM[551] = 32'h05540871,
        RAM[552] = 32'h70840553,
        RAM[553] = 32'h0c727084,
        RAM[554] = 32'h05540871,
        RAM[555] = 32'h70840553,
        RAM[556] = 32'h0cf01252,
        RAM[557] = 32'h718f26c9,
        RAM[558] = 32'h38837227,
        RAM[559] = 32'h95387270,
        RAM[560] = 32'h84055408,
        RAM[561] = 32'h71708405,
        RAM[562] = 32'h530cfc12,
        RAM[563] = 32'h52718326,
        RAM[564] = 32'hed387054,
        RAM[565] = 32'hff8339f7,
        RAM[566] = 32'h3d0d7c70,
        RAM[567] = 32'h525380ca,
        RAM[568] = 32'h3f725490,
        RAM[569] = 32'h08550b0b,
        RAM[570] = 32'h80ce9c56,
        RAM[571] = 32'h81579008,
        RAM[572] = 32'h81055a8b,
        RAM[573] = 32'h3de41159,
        RAM[574] = 32'h538259f4,
        RAM[575] = 32'h13527b88,
        RAM[576] = 32'h11085253,
        RAM[577] = 32'h81833f90,
        RAM[578] = 32'h08307090,
        RAM[579] = 32'h08079f2c,
        RAM[580] = 32'h8a07900c,
        RAM[581] = 32'h538b3d0d,
        RAM[582] = 32'h04ff3d0d,
        RAM[583] = 32'h735280cf,
        RAM[584] = 32'hc00851ff,
        RAM[585] = 32'hb23f833d,
        RAM[586] = 32'h0d04fd3d,
        RAM[587] = 32'h0d757071,
        RAM[588] = 32'h83065355,
        RAM[589] = 32'h5270b838,
        RAM[590] = 32'h71700870,
        RAM[591] = 32'h09f7fbfd,
        RAM[592] = 32'hff120670,
        RAM[593] = 32'hf8848281,
        RAM[594] = 32'h80065151,
        RAM[595] = 32'h5253709d,
        RAM[596] = 32'h38841370,
        RAM[597] = 32'h087009f7,
        RAM[598] = 32'hfbfdff12,
        RAM[599] = 32'h0670f884,
        RAM[600] = 32'h82818006,
        RAM[601] = 32'h51515253,
        RAM[602] = 32'h70802ee5,
        RAM[603] = 32'h38725271,
        RAM[604] = 32'h33517080,
        RAM[605] = 32'h2e8a3881,
        RAM[606] = 32'h12703352,
        RAM[607] = 32'h5270f838,
        RAM[608] = 32'h71743190,
        RAM[609] = 32'h0c853d0d,
        RAM[610] = 32'h04f23d0d,
        RAM[611] = 32'h60628811,
        RAM[612] = 32'h08705757,
        RAM[613] = 32'h5f5a7480,
        RAM[614] = 32'h2e818f38,
        RAM[615] = 32'h8c1a2270,
        RAM[616] = 32'h832a8132,
        RAM[617] = 32'h70810651,
        RAM[618] = 32'h55587386,
        RAM[619] = 32'h38901a08,
        RAM[620] = 32'h91387951,
        RAM[621] = 32'h90a13fff,
        RAM[622] = 32'h54900880,
        RAM[623] = 32'hed388c1a,
        RAM[624] = 32'h22587d08,
        RAM[625] = 32'h57807883,
        RAM[626] = 32'hffff0670,
        RAM[627] = 32'h812a7081,
        RAM[628] = 32'h06515657,
        RAM[629] = 32'h5573752e,
        RAM[630] = 32'h80d73874,
        RAM[631] = 32'h90387608,
        RAM[632] = 32'h84180888,
        RAM[633] = 32'h19595659,
        RAM[634] = 32'h74802ef2,
        RAM[635] = 32'h38745488,
        RAM[636] = 32'h80752784,
        RAM[637] = 32'h38888054,
        RAM[638] = 32'h73537852,
        RAM[639] = 32'h9c1a0851,
        RAM[640] = 32'ha41a0854,
        RAM[641] = 32'h732d800b,
        RAM[642] = 32'h90082582,
        RAM[643] = 32'he6389008,
        RAM[644] = 32'h19759008,
        RAM[645] = 32'h317f8805,
        RAM[646] = 32'h08900831,
        RAM[647] = 32'h70618805,
        RAM[648] = 32'h0c565659,
        RAM[649] = 32'h73ffb438,
        RAM[650] = 32'h80547390,
        RAM[651] = 32'h0c903d0d,
        RAM[652] = 32'h04758132,
        RAM[653] = 32'h70810676,
        RAM[654] = 32'h41515473,
        RAM[655] = 32'h802e81c1,
        RAM[656] = 32'h38749038,
        RAM[657] = 32'h76088418,
        RAM[658] = 32'h08881959,
        RAM[659] = 32'h56597480,
        RAM[660] = 32'h2ef23888,
        RAM[661] = 32'h1a087883,
        RAM[662] = 32'hffff0670,
        RAM[663] = 32'h892a7081,
        RAM[664] = 32'h06515659,
        RAM[665] = 32'h5673802e,
        RAM[666] = 32'h82fa3875,
        RAM[667] = 32'h75278d38,
        RAM[668] = 32'h77872a70,
        RAM[669] = 32'h81065154,
        RAM[670] = 32'h7382b538,
        RAM[671] = 32'h74762783,
        RAM[672] = 32'h38745675,
        RAM[673] = 32'h53785279,
        RAM[674] = 32'h08518582,
        RAM[675] = 32'h3f881a08,
        RAM[676] = 32'h7631881b,
        RAM[677] = 32'h0c790816,
        RAM[678] = 32'h7a0c7456,
        RAM[679] = 32'h75197577,
        RAM[680] = 32'h317f8805,
        RAM[681] = 32'h08783170,
        RAM[682] = 32'h6188050c,
        RAM[683] = 32'h56565973,
        RAM[684] = 32'h802efef4,
        RAM[685] = 32'h388c1a22,
        RAM[686] = 32'h58ff8639,
        RAM[687] = 32'h77785479,
        RAM[688] = 32'h537b5256,
        RAM[689] = 32'h84c83f88,
        RAM[690] = 32'h1a087831,
        RAM[691] = 32'h881b0c79,
        RAM[692] = 32'h08187a0c,
        RAM[693] = 32'h7c76315d,
        RAM[694] = 32'h7c8e3879,
        RAM[695] = 32'h518fdb3f,
        RAM[696] = 32'h9008818f,
        RAM[697] = 32'h3890085f,
        RAM[698] = 32'h75197577,
        RAM[699] = 32'h317f8805,
        RAM[700] = 32'h08783170,
        RAM[701] = 32'h6188050c,
        RAM[702] = 32'h56565973,
        RAM[703] = 32'h802efea8,
        RAM[704] = 32'h38748183,
        RAM[705] = 32'h38760884,
        RAM[706] = 32'h18088819,
        RAM[707] = 32'h59565974,
        RAM[708] = 32'h802ef238,
        RAM[709] = 32'h74538a52,
        RAM[710] = 32'h785182d3,
        RAM[711] = 32'h3f900879,
        RAM[712] = 32'h3181055d,
        RAM[713] = 32'h90088438,
        RAM[714] = 32'h81155d81,
        RAM[715] = 32'h5f7c5874,
        RAM[716] = 32'h7d278338,
        RAM[717] = 32'h7458941a,
        RAM[718] = 32'h08881b08,
        RAM[719] = 32'h11575c80,
        RAM[720] = 32'h7a085c54,
        RAM[721] = 32'h901a087b,
        RAM[722] = 32'h27833881,
        RAM[723] = 32'h54757825,
        RAM[724] = 32'h843873ba,
        RAM[725] = 32'h387b7824,
        RAM[726] = 32'hfee2387b,
        RAM[727] = 32'h5378529c,
        RAM[728] = 32'h1a0851a4,
        RAM[729] = 32'h1a085473,
        RAM[730] = 32'h2d900856,
        RAM[731] = 32'h90088024,
        RAM[732] = 32'hfee2388c,
        RAM[733] = 32'h1a2280c0,
        RAM[734] = 32'h0754738c,
        RAM[735] = 32'h1b23ff54,
        RAM[736] = 32'h73900c90,
        RAM[737] = 32'h3d0d047e,
        RAM[738] = 32'hffa338ff,
        RAM[739] = 32'h87397553,
        RAM[740] = 32'h78527a51,
        RAM[741] = 32'h82f83f79,
        RAM[742] = 32'h08167a0c,
        RAM[743] = 32'h79518e9a,
        RAM[744] = 32'h3f9008cf,
        RAM[745] = 32'h387c7631,
        RAM[746] = 32'h5d7cfebc,
        RAM[747] = 32'h38feac39,
        RAM[748] = 32'h901a087a,
        RAM[749] = 32'h08713176,
        RAM[750] = 32'h1170565a,
        RAM[751] = 32'h575280cf,
        RAM[752] = 32'hc0085184,
        RAM[753] = 32'h8c3f9008,
        RAM[754] = 32'h802effa7,
        RAM[755] = 32'h38900890,
        RAM[756] = 32'h1b0c9008,
        RAM[757] = 32'h167a0c77,
        RAM[758] = 32'h941b0c74,
        RAM[759] = 32'h881b0c74,
        RAM[760] = 32'h56fd9939,
        RAM[761] = 32'h79085890,
        RAM[762] = 32'h1a087827,
        RAM[763] = 32'h83388154,
        RAM[764] = 32'h75752784,
        RAM[765] = 32'h3873b338,
        RAM[766] = 32'h941a0856,
        RAM[767] = 32'h75752680,
        RAM[768] = 32'hd3387553,
        RAM[769] = 32'h78529c1a,
        RAM[770] = 32'h0851a41a,
        RAM[771] = 32'h0854732d,
        RAM[772] = 32'h90085690,
        RAM[773] = 32'h088024fd,
        RAM[774] = 32'h83388c1a,
        RAM[775] = 32'h2280c007,
        RAM[776] = 32'h54738c1b,
        RAM[777] = 32'h23ff54fe,
        RAM[778] = 32'hd7397553,
        RAM[779] = 32'h78527751,
        RAM[780] = 32'h81dc3f79,
        RAM[781] = 32'h08167a0c,
        RAM[782] = 32'h79518cfe,
        RAM[783] = 32'h3f900880,
        RAM[784] = 32'h2efcd938,
        RAM[785] = 32'h8c1a2280,
        RAM[786] = 32'hc0075473,
        RAM[787] = 32'h8c1b23ff,
        RAM[788] = 32'h54fead39,
        RAM[789] = 32'h74755479,
        RAM[790] = 32'h53785256,
        RAM[791] = 32'h81b03f88,
        RAM[792] = 32'h1a087531,
        RAM[793] = 32'h881b0c79,
        RAM[794] = 32'h08157a0c,
        RAM[795] = 32'hfcae39fa,
        RAM[796] = 32'h3d0d7a79,
        RAM[797] = 32'h028805a7,
        RAM[798] = 32'h05335652,
        RAM[799] = 32'h53837327,
        RAM[800] = 32'h8a387083,
        RAM[801] = 32'h06527180,
        RAM[802] = 32'h2ea838ff,
        RAM[803] = 32'h135372ff,
        RAM[804] = 32'h2e973870,
        RAM[805] = 32'h33527372,
        RAM[806] = 32'h2e913881,
        RAM[807] = 32'h11ff1454,
        RAM[808] = 32'h5172ff2e,
        RAM[809] = 32'h098106eb,
        RAM[810] = 32'h38805170,
        RAM[811] = 32'h900c883d,
        RAM[812] = 32'h0d047072,
        RAM[813] = 32'h57558351,
        RAM[814] = 32'h75828029,
        RAM[815] = 32'h14ff1252,
        RAM[816] = 32'h56708025,
        RAM[817] = 32'hf3388373,
        RAM[818] = 32'h27bf3874,
        RAM[819] = 32'h08763270,
        RAM[820] = 32'h09f7fbfd,
        RAM[821] = 32'hff120670,
        RAM[822] = 32'hf8848281,
        RAM[823] = 32'h80065151,
        RAM[824] = 32'h5170802e,
        RAM[825] = 32'h99387451,
        RAM[826] = 32'h80527033,
        RAM[827] = 32'h5773772e,
        RAM[828] = 32'hffb93881,
        RAM[829] = 32'h11811353,
        RAM[830] = 32'h51837227,
        RAM[831] = 32'hed38fc13,
        RAM[832] = 32'h84165653,
        RAM[833] = 32'h728326c3,
        RAM[834] = 32'h387451fe,
        RAM[835] = 32'hfe39fa3d,
        RAM[836] = 32'h0d787a7c,
        RAM[837] = 32'h72727257,
        RAM[838] = 32'h57575956,
        RAM[839] = 32'h56747627,
        RAM[840] = 32'hb2387615,
        RAM[841] = 32'h51757127,
        RAM[842] = 32'haa387077,
        RAM[843] = 32'h17ff1454,
        RAM[844] = 32'h555371ff,
        RAM[845] = 32'h2e9638ff,
        RAM[846] = 32'h14ff1454,
        RAM[847] = 32'h54723374,
        RAM[848] = 32'h34ff1252,
        RAM[849] = 32'h71ff2e09,
        RAM[850] = 32'h8106ec38,
        RAM[851] = 32'h75900c88,
        RAM[852] = 32'h3d0d0476,
        RAM[853] = 32'h8f269738,
        RAM[854] = 32'hff125271,
        RAM[855] = 32'hff2eed38,
        RAM[856] = 32'h72708105,
        RAM[857] = 32'h54337470,
        RAM[858] = 32'h81055634,
        RAM[859] = 32'heb397476,
        RAM[860] = 32'h07830651,
        RAM[861] = 32'h70e23875,
        RAM[862] = 32'h75545172,
        RAM[863] = 32'h70840554,
        RAM[864] = 32'h08717084,
        RAM[865] = 32'h05530c72,
        RAM[866] = 32'h70840554,
        RAM[867] = 32'h08717084,
        RAM[868] = 32'h05530c72,
        RAM[869] = 32'h70840554,
        RAM[870] = 32'h08717084,
        RAM[871] = 32'h05530c72,
        RAM[872] = 32'h70840554,
        RAM[873] = 32'h08717084,
        RAM[874] = 32'h05530cf0,
        RAM[875] = 32'h1252718f,
        RAM[876] = 32'h26c93883,
        RAM[877] = 32'h72279538,
        RAM[878] = 32'h72708405,
        RAM[879] = 32'h54087170,
        RAM[880] = 32'h8405530c,
        RAM[881] = 32'hfc125271,
        RAM[882] = 32'h8326ed38,
        RAM[883] = 32'h7054ff88,
        RAM[884] = 32'h39ef3d0d,
        RAM[885] = 32'h63656740,
        RAM[886] = 32'h5d427b80,
        RAM[887] = 32'h2e84fa38,
        RAM[888] = 32'h6151a5b4,
        RAM[889] = 32'h3ff81c70,
        RAM[890] = 32'h84120870,
        RAM[891] = 32'hfc067062,
        RAM[892] = 32'h8b0570f8,
        RAM[893] = 32'h06415945,
        RAM[894] = 32'h5b5c4157,
        RAM[895] = 32'h96742782,
        RAM[896] = 32'hc338807b,
        RAM[897] = 32'h247e7c26,
        RAM[898] = 32'h07598054,
        RAM[899] = 32'h78742e09,
        RAM[900] = 32'h810682a9,
        RAM[901] = 32'h38777b25,
        RAM[902] = 32'h81fc3877,
        RAM[903] = 32'h1780d6fc,
        RAM[904] = 32'h0b880508,
        RAM[905] = 32'h5e567c76,
        RAM[906] = 32'h2e84bd38,
        RAM[907] = 32'h84160870,
        RAM[908] = 32'hfe061784,
        RAM[909] = 32'h11088106,
        RAM[910] = 32'h51555573,
        RAM[911] = 32'h828b3874,
        RAM[912] = 32'hfc06597c,
        RAM[913] = 32'h762e84dd,
        RAM[914] = 32'h3877195f,
        RAM[915] = 32'h7e7b2581,
        RAM[916] = 32'hfd387981,
        RAM[917] = 32'h06547382,
        RAM[918] = 32'hbf387677,
        RAM[919] = 32'h08318411,
        RAM[920] = 32'h08fc0656,
        RAM[921] = 32'h5a75802e,
        RAM[922] = 32'h91387c76,
        RAM[923] = 32'h2e84ea38,
        RAM[924] = 32'h74191859,
        RAM[925] = 32'h787b2584,
        RAM[926] = 32'h89387980,
        RAM[927] = 32'h2e829938,
        RAM[928] = 32'h7715567a,
        RAM[929] = 32'h76248290,
        RAM[930] = 32'h388c1a08,
        RAM[931] = 32'h881b0871,
        RAM[932] = 32'h8c120c88,
        RAM[933] = 32'h120c5579,
        RAM[934] = 32'h76595788,
        RAM[935] = 32'h1761fc05,
        RAM[936] = 32'h575975a4,
        RAM[937] = 32'h2685ef38,
        RAM[938] = 32'h7b795555,
        RAM[939] = 32'h93762780,
        RAM[940] = 32'hc9387b70,
        RAM[941] = 32'h84055d08,
        RAM[942] = 32'h7c56790c,
        RAM[943] = 32'h74708405,
        RAM[944] = 32'h56088c18,
        RAM[945] = 32'h0c901754,
        RAM[946] = 32'h9b7627ae,
        RAM[947] = 32'h38747084,
        RAM[948] = 32'h05560874,
        RAM[949] = 32'h0c747084,
        RAM[950] = 32'h05560894,
        RAM[951] = 32'h180c9817,
        RAM[952] = 32'h54a37627,
        RAM[953] = 32'h95387470,
        RAM[954] = 32'h84055608,
        RAM[955] = 32'h740c7470,
        RAM[956] = 32'h84055608,
        RAM[957] = 32'h9c180ca0,
        RAM[958] = 32'h17547470,
        RAM[959] = 32'h84055608,
        RAM[960] = 32'h74708405,
        RAM[961] = 32'h560c7470,
        RAM[962] = 32'h84055608,
        RAM[963] = 32'h74708405,
        RAM[964] = 32'h560c7408,
        RAM[965] = 32'h740c777b,
        RAM[966] = 32'h3156758f,
        RAM[967] = 32'h2680c938,
        RAM[968] = 32'h84170881,
        RAM[969] = 32'h06780784,
        RAM[970] = 32'h180c7717,
        RAM[971] = 32'h84110881,
        RAM[972] = 32'h0784120c,
        RAM[973] = 32'h546151a2,
        RAM[974] = 32'he03f8817,
        RAM[975] = 32'h5473900c,
        RAM[976] = 32'h933d0d04,
        RAM[977] = 32'h905bfdba,
        RAM[978] = 32'h397856fe,
        RAM[979] = 32'h85398c16,
        RAM[980] = 32'h08881708,
        RAM[981] = 32'h718c120c,
        RAM[982] = 32'h88120c55,
        RAM[983] = 32'h7e707c31,
        RAM[984] = 32'h57588f76,
        RAM[985] = 32'h27ffb938,
        RAM[986] = 32'h7a178418,
        RAM[987] = 32'h0881067c,
        RAM[988] = 32'h0784190c,
        RAM[989] = 32'h76810784,
        RAM[990] = 32'h120c7611,
        RAM[991] = 32'h84110881,
        RAM[992] = 32'h0784120c,
        RAM[993] = 32'h55880552,
        RAM[994] = 32'h61518cf6,
        RAM[995] = 32'h3f6151a2,
        RAM[996] = 32'h883f8817,
        RAM[997] = 32'h54ffa639,
        RAM[998] = 32'h7d526151,
        RAM[999] = 32'h94f53f90,
        RAM[1000] = 32'h08599008,
        RAM[1001] = 32'h802e81a3,
        RAM[1002] = 32'h389008f8,
        RAM[1003] = 32'h05608405,
        RAM[1004] = 32'h08fe0661,
        RAM[1005] = 32'h05555776,
        RAM[1006] = 32'h742e83e6,
        RAM[1007] = 32'h38fc1856,
        RAM[1008] = 32'h75a42681,
        RAM[1009] = 32'haa387b90,
        RAM[1010] = 32'h08555593,
        RAM[1011] = 32'h762780d8,
        RAM[1012] = 32'h38747084,
        RAM[1013] = 32'h05560890,
        RAM[1014] = 32'h08708405,
        RAM[1015] = 32'h900c0c90,
        RAM[1016] = 32'h08757084,
        RAM[1017] = 32'h05570871,
        RAM[1018] = 32'h70840553,
        RAM[1019] = 32'h0c549b76,
        RAM[1020] = 32'h27b63874,
        RAM[1021] = 32'h70840556,
        RAM[1022] = 32'h08747084,
        RAM[1023] = 32'h05560c74,
        RAM[1024] = 32'h70840556,
        RAM[1025] = 32'h08747084,
        RAM[1026] = 32'h05560ca3,
        RAM[1027] = 32'h76279938,
        RAM[1028] = 32'h74708405,
        RAM[1029] = 32'h56087470,
        RAM[1030] = 32'h8405560c,
        RAM[1031] = 32'h74708405,
        RAM[1032] = 32'h56087470,
        RAM[1033] = 32'h8405560c,
        RAM[1034] = 32'h74708405,
        RAM[1035] = 32'h56087470,
        RAM[1036] = 32'h8405560c,
        RAM[1037] = 32'h74708405,
        RAM[1038] = 32'h56087470,
        RAM[1039] = 32'h8405560c,
        RAM[1040] = 32'h7408740c,
        RAM[1041] = 32'h7b526151,
        RAM[1042] = 32'h8bb83f61,
        RAM[1043] = 32'h51a0ca3f,
        RAM[1044] = 32'h78547390,
        RAM[1045] = 32'h0c933d0d,
        RAM[1046] = 32'h047d5261,
        RAM[1047] = 32'h5193b43f,
        RAM[1048] = 32'h9008900c,
        RAM[1049] = 32'h933d0d04,
        RAM[1050] = 32'h84160855,
        RAM[1051] = 32'hfbd13975,
        RAM[1052] = 32'h537b5290,
        RAM[1053] = 32'h0851efc6,
        RAM[1054] = 32'h3f7b5261,
        RAM[1055] = 32'h518b833f,
        RAM[1056] = 32'hca398c16,
        RAM[1057] = 32'h08881708,
        RAM[1058] = 32'h718c120c,
        RAM[1059] = 32'h88120c55,
        RAM[1060] = 32'h8c1a0888,
        RAM[1061] = 32'h1b08718c,
        RAM[1062] = 32'h120c8812,
        RAM[1063] = 32'h0c557979,
        RAM[1064] = 32'h5957fbf7,
        RAM[1065] = 32'h39771990,
        RAM[1066] = 32'h1c555573,
        RAM[1067] = 32'h7524fba2,
        RAM[1068] = 32'h387a1770,
        RAM[1069] = 32'h80d6fc0b,
        RAM[1070] = 32'h88050c75,
        RAM[1071] = 32'h7c318107,
        RAM[1072] = 32'h84120c5d,
        RAM[1073] = 32'h84170881,
        RAM[1074] = 32'h067b0784,
        RAM[1075] = 32'h180c6151,
        RAM[1076] = 32'h9fc73f88,
        RAM[1077] = 32'h1754fce5,
        RAM[1078] = 32'h39741918,
        RAM[1079] = 32'h901c555d,
        RAM[1080] = 32'h737d24fb,
        RAM[1081] = 32'h95388c1a,
        RAM[1082] = 32'h08881b08,
        RAM[1083] = 32'h718c120c,
        RAM[1084] = 32'h88120c55,
        RAM[1085] = 32'h881a61fc,
        RAM[1086] = 32'h05575975,
        RAM[1087] = 32'ha42681ae,
        RAM[1088] = 32'h387b7955,
        RAM[1089] = 32'h55937627,
        RAM[1090] = 32'h80c9387b,
        RAM[1091] = 32'h7084055d,
        RAM[1092] = 32'h087c5679,
        RAM[1093] = 32'h0c747084,
        RAM[1094] = 32'h0556088c,
        RAM[1095] = 32'h1b0c901a,
        RAM[1096] = 32'h549b7627,
        RAM[1097] = 32'hae387470,
        RAM[1098] = 32'h84055608,
        RAM[1099] = 32'h740c7470,
        RAM[1100] = 32'h84055608,
        RAM[1101] = 32'h941b0c98,
        RAM[1102] = 32'h1a54a376,
        RAM[1103] = 32'h27953874,
        RAM[1104] = 32'h70840556,
        RAM[1105] = 32'h08740c74,
        RAM[1106] = 32'h70840556,
        RAM[1107] = 32'h089c1b0c,
        RAM[1108] = 32'ha01a5474,
        RAM[1109] = 32'h70840556,
        RAM[1110] = 32'h08747084,
        RAM[1111] = 32'h05560c74,
        RAM[1112] = 32'h70840556,
        RAM[1113] = 32'h08747084,
        RAM[1114] = 32'h05560c74,
        RAM[1115] = 32'h08740c7a,
        RAM[1116] = 32'h1a7080d6,
        RAM[1117] = 32'hfc0b8805,
        RAM[1118] = 32'h0c7d7c31,
        RAM[1119] = 32'h81078412,
        RAM[1120] = 32'h0c54841a,
        RAM[1121] = 32'h0881067b,
        RAM[1122] = 32'h07841b0c,
        RAM[1123] = 32'h61519e89,
        RAM[1124] = 32'h3f7854fd,
        RAM[1125] = 32'hbd397553,
        RAM[1126] = 32'h7b527851,
        RAM[1127] = 32'heda03ffa,
        RAM[1128] = 32'hf5398417,
        RAM[1129] = 32'h08fc0618,
        RAM[1130] = 32'h605858fa,
        RAM[1131] = 32'he9397553,
        RAM[1132] = 32'h7b527851,
        RAM[1133] = 32'hed883f7a,
        RAM[1134] = 32'h1a7080d6,
        RAM[1135] = 32'hfc0b8805,
        RAM[1136] = 32'h0c7d7c31,
        RAM[1137] = 32'h81078412,
        RAM[1138] = 32'h0c54841a,
        RAM[1139] = 32'h0881067b,
        RAM[1140] = 32'h07841b0c,
        RAM[1141] = 32'hffb639fa,
        RAM[1142] = 32'h3d0d7880,
        RAM[1143] = 32'hcfc00854,
        RAM[1144] = 32'h55b81308,
        RAM[1145] = 32'h802e81b5,
        RAM[1146] = 32'h388c1522,
        RAM[1147] = 32'h7083ffff,
        RAM[1148] = 32'h0670832a,
        RAM[1149] = 32'h81327081,
        RAM[1150] = 32'h06515555,
        RAM[1151] = 32'h5672802e,
        RAM[1152] = 32'h80dc3873,
        RAM[1153] = 32'h842a8132,
        RAM[1154] = 32'h810657ff,
        RAM[1155] = 32'h537680f6,
        RAM[1156] = 32'h3873822a,
        RAM[1157] = 32'h70810651,
        RAM[1158] = 32'h5372802e,
        RAM[1159] = 32'hb938b015,
        RAM[1160] = 32'h08547380,
        RAM[1161] = 32'h2e9c3880,
        RAM[1162] = 32'hc0155373,
        RAM[1163] = 32'h732e8f38,
        RAM[1164] = 32'h735280cf,
        RAM[1165] = 32'hc0085187,
        RAM[1166] = 32'hc93f8c15,
        RAM[1167] = 32'h225676b0,
        RAM[1168] = 32'h160c75db,
        RAM[1169] = 32'h0653728c,
        RAM[1170] = 32'h1623800b,
        RAM[1171] = 32'h84160c90,
        RAM[1172] = 32'h1508750c,
        RAM[1173] = 32'h72567588,
        RAM[1174] = 32'h0753728c,
        RAM[1175] = 32'h16239015,
        RAM[1176] = 32'h08802e80,
        RAM[1177] = 32'hc0388c15,
        RAM[1178] = 32'h22708106,
        RAM[1179] = 32'h5553739d,
        RAM[1180] = 32'h3872812a,
        RAM[1181] = 32'h70810651,
        RAM[1182] = 32'h53728538,
        RAM[1183] = 32'h94150854,
        RAM[1184] = 32'h7388160c,
        RAM[1185] = 32'h80537290,
        RAM[1186] = 32'h0c883d0d,
        RAM[1187] = 32'h04800b88,
        RAM[1188] = 32'h160c9415,
        RAM[1189] = 32'h08309816,
        RAM[1190] = 32'h0c8053ea,
        RAM[1191] = 32'h39725182,
        RAM[1192] = 32'hfb3ffec5,
        RAM[1193] = 32'h3974518c,
        RAM[1194] = 32'he83f8c15,
        RAM[1195] = 32'h22708106,
        RAM[1196] = 32'h55537380,
        RAM[1197] = 32'h2effba38,
        RAM[1198] = 32'hd439f83d,
        RAM[1199] = 32'h0d7a5877,
        RAM[1200] = 32'h802e8199,
        RAM[1201] = 32'h3880cfc0,
        RAM[1202] = 32'h0854b814,
        RAM[1203] = 32'h08802e80,
        RAM[1204] = 32'hed388c18,
        RAM[1205] = 32'h2270902b,
        RAM[1206] = 32'h70902c70,
        RAM[1207] = 32'h832a8132,
        RAM[1208] = 32'h81065c51,
        RAM[1209] = 32'h57547880,
        RAM[1210] = 32'hcd389018,
        RAM[1211] = 32'h08577680,
        RAM[1212] = 32'h2e80c338,
        RAM[1213] = 32'h77087731,
        RAM[1214] = 32'h77790c76,
        RAM[1215] = 32'h83067a58,
        RAM[1216] = 32'h55557385,
        RAM[1217] = 32'h38941808,
        RAM[1218] = 32'h56758819,
        RAM[1219] = 32'h0c807525,
        RAM[1220] = 32'ha5387453,
        RAM[1221] = 32'h76529c18,
        RAM[1222] = 32'h0851a418,
        RAM[1223] = 32'h0854732d,
        RAM[1224] = 32'h800b9008,
        RAM[1225] = 32'h2580c938,
        RAM[1226] = 32'h90081775,
        RAM[1227] = 32'h90083156,
        RAM[1228] = 32'h57748024,
        RAM[1229] = 32'hdd38800b,
        RAM[1230] = 32'h900c8a3d,
        RAM[1231] = 32'h0d047351,
        RAM[1232] = 32'h81da3f8c,
        RAM[1233] = 32'h18227090,
        RAM[1234] = 32'h2b70902c,
        RAM[1235] = 32'h70832a81,
        RAM[1236] = 32'h3281065c,
        RAM[1237] = 32'h51575478,
        RAM[1238] = 32'hdd38ff8e,
        RAM[1239] = 32'h39a5b652,
        RAM[1240] = 32'h80cfc008,
        RAM[1241] = 32'h5189f13f,
        RAM[1242] = 32'h9008900c,
        RAM[1243] = 32'h8a3d0d04,
        RAM[1244] = 32'h8c182280,
        RAM[1245] = 32'hc0075473,
        RAM[1246] = 32'h8c1923ff,
        RAM[1247] = 32'h0b900c8a,
        RAM[1248] = 32'h3d0d0480,
        RAM[1249] = 32'h3d0d7251,
        RAM[1250] = 32'h80710c80,
        RAM[1251] = 32'h0b84120c,
        RAM[1252] = 32'h800b8812,
        RAM[1253] = 32'h0c028e05,
        RAM[1254] = 32'h228c1223,
        RAM[1255] = 32'h02920522,
        RAM[1256] = 32'h8e122380,
        RAM[1257] = 32'h0b90120c,
        RAM[1258] = 32'h800b9412,
        RAM[1259] = 32'h0c800b98,
        RAM[1260] = 32'h120c709c,
        RAM[1261] = 32'h120c80c1,
        RAM[1262] = 32'hca0ba012,
        RAM[1263] = 32'h0c80c296,
        RAM[1264] = 32'h0ba4120c,
        RAM[1265] = 32'h80c3920b,
        RAM[1266] = 32'ha8120c80,
        RAM[1267] = 32'hc3e30bac,
        RAM[1268] = 32'h120c823d,
        RAM[1269] = 32'h0d04fa3d,
        RAM[1270] = 32'h0d797080,
        RAM[1271] = 32'hdc298c11,
        RAM[1272] = 32'h547a5356,
        RAM[1273] = 32'h578cac3f,
        RAM[1274] = 32'h90089008,
        RAM[1275] = 32'h55569008,
        RAM[1276] = 32'h802ea238,
        RAM[1277] = 32'h90088c05,
        RAM[1278] = 32'h54800b90,
        RAM[1279] = 32'h080c7690,
        RAM[1280] = 32'h0884050c,
        RAM[1281] = 32'h73900888,
        RAM[1282] = 32'h050c7453,
        RAM[1283] = 32'h80527351,
        RAM[1284] = 32'h97f73f75,
        RAM[1285] = 32'h5473900c,
        RAM[1286] = 32'h883d0d04,
        RAM[1287] = 32'hfc3d0d76,
        RAM[1288] = 32'haaab0bbc,
        RAM[1289] = 32'h120c5581,
        RAM[1290] = 32'h0bb8160c,
        RAM[1291] = 32'h800b84dc,
        RAM[1292] = 32'h160c830b,
        RAM[1293] = 32'h84e0160c,
        RAM[1294] = 32'h84e81584,
        RAM[1295] = 32'he4160c74,
        RAM[1296] = 32'h54805384,
        RAM[1297] = 32'h52841508,
        RAM[1298] = 32'h51feb83f,
        RAM[1299] = 32'h74548153,
        RAM[1300] = 32'h89528815,
        RAM[1301] = 32'h0851feab,
        RAM[1302] = 32'h3f745482,
        RAM[1303] = 32'h538a528c,
        RAM[1304] = 32'h150851fe,
        RAM[1305] = 32'h9e3f863d,
        RAM[1306] = 32'h0d04f93d,
        RAM[1307] = 32'h0d7980cf,
        RAM[1308] = 32'hc0085457,
        RAM[1309] = 32'hb8130880,
        RAM[1310] = 32'h2e80c838,
        RAM[1311] = 32'h84dc1356,
        RAM[1312] = 32'h88160884,
        RAM[1313] = 32'h1708ff05,
        RAM[1314] = 32'h55558074,
        RAM[1315] = 32'h249f388c,
        RAM[1316] = 32'h15227090,
        RAM[1317] = 32'h2b70902c,
        RAM[1318] = 32'h51545872,
        RAM[1319] = 32'h802e80ca,
        RAM[1320] = 32'h3880dc15,
        RAM[1321] = 32'hff155555,
        RAM[1322] = 32'h738025e3,
        RAM[1323] = 32'h38750853,
        RAM[1324] = 32'h72802e9f,
        RAM[1325] = 32'h38725688,
        RAM[1326] = 32'h16088417,
        RAM[1327] = 32'h08ff0555,
        RAM[1328] = 32'h55c83972,
        RAM[1329] = 32'h51fed53f,
        RAM[1330] = 32'h80cfc008,
        RAM[1331] = 32'h84dc0556,
        RAM[1332] = 32'hffae3984,
        RAM[1333] = 32'h527651fd,
        RAM[1334] = 32'hfd3f9008,
        RAM[1335] = 32'h760c9008,
        RAM[1336] = 32'h802e80c0,
        RAM[1337] = 32'h38900856,
        RAM[1338] = 32'hce39810b,
        RAM[1339] = 32'h8c162372,
        RAM[1340] = 32'h750c7288,
        RAM[1341] = 32'h160c7284,
        RAM[1342] = 32'h160c7290,
        RAM[1343] = 32'h160c7294,
        RAM[1344] = 32'h160c7298,
        RAM[1345] = 32'h160cff0b,
        RAM[1346] = 32'h8e162372,
        RAM[1347] = 32'hb0160c72,
        RAM[1348] = 32'hb4160c72,
        RAM[1349] = 32'h80c4160c,
        RAM[1350] = 32'h7280c816,
        RAM[1351] = 32'h0c74900c,
        RAM[1352] = 32'h893d0d04,
        RAM[1353] = 32'h8c770c80,
        RAM[1354] = 32'h0b900c89,
        RAM[1355] = 32'h3d0d04ff,
        RAM[1356] = 32'h3d0da5b6,
        RAM[1357] = 32'h52735186,
        RAM[1358] = 32'h9f3f833d,
        RAM[1359] = 32'h0d04803d,
        RAM[1360] = 32'h0d80cfc0,
        RAM[1361] = 32'h0851e83f,
        RAM[1362] = 32'h823d0d04,
        RAM[1363] = 32'hfb3d0d77,
        RAM[1364] = 32'h70525696,
        RAM[1365] = 32'hc33f80d6,
        RAM[1366] = 32'hfc0b8805,
        RAM[1367] = 32'h08841108,
        RAM[1368] = 32'hfc06707b,
        RAM[1369] = 32'h319fef05,
        RAM[1370] = 32'he08006e0,
        RAM[1371] = 32'h80055656,
        RAM[1372] = 32'h53a08074,
        RAM[1373] = 32'h24943880,
        RAM[1374] = 32'h52755196,
        RAM[1375] = 32'h9d3f80d7,
        RAM[1376] = 32'h84081553,
        RAM[1377] = 32'h7290082e,
        RAM[1378] = 32'h8f387551,
        RAM[1379] = 32'h968b3f80,
        RAM[1380] = 32'h5372900c,
        RAM[1381] = 32'h873d0d04,
        RAM[1382] = 32'h73305275,
        RAM[1383] = 32'h5195fb3f,
        RAM[1384] = 32'h9008ff2e,
        RAM[1385] = 32'ha83880d6,
        RAM[1386] = 32'hfc0b8805,
        RAM[1387] = 32'h08757531,
        RAM[1388] = 32'h81078412,
        RAM[1389] = 32'h0c5380d6,
        RAM[1390] = 32'hc0087431,
        RAM[1391] = 32'h80d6c00c,
        RAM[1392] = 32'h755195d5,
        RAM[1393] = 32'h3f810b90,
        RAM[1394] = 32'h0c873d0d,
        RAM[1395] = 32'h04805275,
        RAM[1396] = 32'h5195c73f,
        RAM[1397] = 32'h80d6fc0b,
        RAM[1398] = 32'h88050890,
        RAM[1399] = 32'h08713156,
        RAM[1400] = 32'h538f7525,
        RAM[1401] = 32'hffa43890,
        RAM[1402] = 32'h0880d6f0,
        RAM[1403] = 32'h083180d6,
        RAM[1404] = 32'hc00c7481,
        RAM[1405] = 32'h0784140c,
        RAM[1406] = 32'h7551959d,
        RAM[1407] = 32'h3f8053ff,
        RAM[1408] = 32'h9039f63d,
        RAM[1409] = 32'h0d7c7e54,
        RAM[1410] = 32'h5b72802e,
        RAM[1411] = 32'h8283387a,
        RAM[1412] = 32'h5195853f,
        RAM[1413] = 32'hf8138411,
        RAM[1414] = 32'h0870fe06,
        RAM[1415] = 32'h70138411,
        RAM[1416] = 32'h08fc065d,
        RAM[1417] = 32'h58595458,
        RAM[1418] = 32'h80d78408,
        RAM[1419] = 32'h752e82de,
        RAM[1420] = 32'h38788416,
        RAM[1421] = 32'h0c807381,
        RAM[1422] = 32'h06545a72,
        RAM[1423] = 32'h7a2e81d5,
        RAM[1424] = 32'h38781584,
        RAM[1425] = 32'h11088106,
        RAM[1426] = 32'h515372a0,
        RAM[1427] = 32'h38781757,
        RAM[1428] = 32'h7981e638,
        RAM[1429] = 32'h88150853,
        RAM[1430] = 32'h7280d784,
        RAM[1431] = 32'h2e82f938,
        RAM[1432] = 32'h8c150870,
        RAM[1433] = 32'h8c150c73,
        RAM[1434] = 32'h88120c56,
        RAM[1435] = 32'h76810784,
        RAM[1436] = 32'h190c7618,
        RAM[1437] = 32'h77710c53,
        RAM[1438] = 32'h79819138,
        RAM[1439] = 32'h83ff7727,
        RAM[1440] = 32'h81c83876,
        RAM[1441] = 32'h892a7783,
        RAM[1442] = 32'h2a565372,
        RAM[1443] = 32'h802ebf38,
        RAM[1444] = 32'h76862ab8,
        RAM[1445] = 32'h05558473,
        RAM[1446] = 32'h27b43880,
        RAM[1447] = 32'hdb135594,
        RAM[1448] = 32'h7327ab38,
        RAM[1449] = 32'h768c2a80,
        RAM[1450] = 32'hee055580,
        RAM[1451] = 32'hd473279e,
        RAM[1452] = 32'h38768f2a,
        RAM[1453] = 32'h80f70555,
        RAM[1454] = 32'h82d47327,
        RAM[1455] = 32'h91387692,
        RAM[1456] = 32'h2a80fc05,
        RAM[1457] = 32'h558ad473,
        RAM[1458] = 32'h27843880,
        RAM[1459] = 32'hfe557410,
        RAM[1460] = 32'h101080d6,
        RAM[1461] = 32'hfc058811,
        RAM[1462] = 32'h08555673,
        RAM[1463] = 32'h762e82b3,
        RAM[1464] = 32'h38841408,
        RAM[1465] = 32'hfc065376,
        RAM[1466] = 32'h73278d38,
        RAM[1467] = 32'h88140854,
        RAM[1468] = 32'h73762e09,
        RAM[1469] = 32'h8106ea38,
        RAM[1470] = 32'h8c140870,
        RAM[1471] = 32'h8c1a0c74,
        RAM[1472] = 32'h881a0c78,
        RAM[1473] = 32'h88120c56,
        RAM[1474] = 32'h778c150c,
        RAM[1475] = 32'h7a519389,
        RAM[1476] = 32'h3f8c3d0d,
        RAM[1477] = 32'h04770878,
        RAM[1478] = 32'h71315977,
        RAM[1479] = 32'h05881908,
        RAM[1480] = 32'h54577280,
        RAM[1481] = 32'hd7842e80,
        RAM[1482] = 32'he0388c18,
        RAM[1483] = 32'h08708c15,
        RAM[1484] = 32'h0c738812,
        RAM[1485] = 32'h0c56fe89,
        RAM[1486] = 32'h39881508,
        RAM[1487] = 32'h8c160870,
        RAM[1488] = 32'h8c130c57,
        RAM[1489] = 32'h88170cfe,
        RAM[1490] = 32'ha3397683,
        RAM[1491] = 32'h2a705455,
        RAM[1492] = 32'h80752481,
        RAM[1493] = 32'h98387282,
        RAM[1494] = 32'h2c81712b,
        RAM[1495] = 32'h80d78008,
        RAM[1496] = 32'h0780d6fc,
        RAM[1497] = 32'h0b84050c,
        RAM[1498] = 32'h53741010,
        RAM[1499] = 32'h1080d6fc,
        RAM[1500] = 32'h05881108,
        RAM[1501] = 32'h5556758c,
        RAM[1502] = 32'h190c7388,
        RAM[1503] = 32'h190c7788,
        RAM[1504] = 32'h170c778c,
        RAM[1505] = 32'h150cff84,
        RAM[1506] = 32'h39815afd,
        RAM[1507] = 32'hb4397817,
        RAM[1508] = 32'h73810654,
        RAM[1509] = 32'h57729838,
        RAM[1510] = 32'h77087871,
        RAM[1511] = 32'h31597705,
        RAM[1512] = 32'h8c190888,
        RAM[1513] = 32'h1a08718c,
        RAM[1514] = 32'h120c8812,
        RAM[1515] = 32'h0c575776,
        RAM[1516] = 32'h81078419,
        RAM[1517] = 32'h0c7780d6,
        RAM[1518] = 32'hfc0b8805,
        RAM[1519] = 32'h0c80d6f8,
        RAM[1520] = 32'h087726fe,
        RAM[1521] = 32'hc73880d6,
        RAM[1522] = 32'hf408527a,
        RAM[1523] = 32'h51fafd3f,
        RAM[1524] = 32'h7a5191c5,
        RAM[1525] = 32'h3ffeba39,
        RAM[1526] = 32'h81788c15,
        RAM[1527] = 32'h0c788815,
        RAM[1528] = 32'h0c738c1a,
        RAM[1529] = 32'h0c73881a,
        RAM[1530] = 32'h0c5afd80,
        RAM[1531] = 32'h39831570,
        RAM[1532] = 32'h822c8171,
        RAM[1533] = 32'h2b80d780,
        RAM[1534] = 32'h080780d6,
        RAM[1535] = 32'hfc0b8405,
        RAM[1536] = 32'h0c515374,
        RAM[1537] = 32'h10101080,
        RAM[1538] = 32'hd6fc0588,
        RAM[1539] = 32'h11085556,
        RAM[1540] = 32'hfee43974,
        RAM[1541] = 32'h53807524,
        RAM[1542] = 32'ha7387282,
        RAM[1543] = 32'h2c81712b,
        RAM[1544] = 32'h80d78008,
        RAM[1545] = 32'h0780d6fc,
        RAM[1546] = 32'h0b84050c,
        RAM[1547] = 32'h53758c19,
        RAM[1548] = 32'h0c738819,
        RAM[1549] = 32'h0c778817,
        RAM[1550] = 32'h0c778c15,
        RAM[1551] = 32'h0cfdcd39,
        RAM[1552] = 32'h83157082,
        RAM[1553] = 32'h2c81712b,
        RAM[1554] = 32'h80d78008,
        RAM[1555] = 32'h0780d6fc,
        RAM[1556] = 32'h0b84050c,
        RAM[1557] = 32'h5153d639,
        RAM[1558] = 32'hf93d0d79,
        RAM[1559] = 32'h7b585380,
        RAM[1560] = 32'h0b80cfc0,
        RAM[1561] = 32'h08535672,
        RAM[1562] = 32'h722e80c0,
        RAM[1563] = 32'h3884dc13,
        RAM[1564] = 32'h5574762e,
        RAM[1565] = 32'hb7388815,
        RAM[1566] = 32'h08841608,
        RAM[1567] = 32'hff055454,
        RAM[1568] = 32'h8073249d,
        RAM[1569] = 32'h388c1422,
        RAM[1570] = 32'h70902b70,
        RAM[1571] = 32'h902c5153,
        RAM[1572] = 32'h587180d8,
        RAM[1573] = 32'h3880dc14,
        RAM[1574] = 32'hff145454,
        RAM[1575] = 32'h728025e5,
        RAM[1576] = 32'h38740855,
        RAM[1577] = 32'h74d03880,
        RAM[1578] = 32'hcfc00852,
        RAM[1579] = 32'h84dc1255,
        RAM[1580] = 32'h74802eb1,
        RAM[1581] = 32'h38881508,
        RAM[1582] = 32'h841608ff,
        RAM[1583] = 32'h05545480,
        RAM[1584] = 32'h73249c38,
        RAM[1585] = 32'h8c142270,
        RAM[1586] = 32'h902b7090,
        RAM[1587] = 32'h2c515358,
        RAM[1588] = 32'h71ad3880,
        RAM[1589] = 32'hdc14ff14,
        RAM[1590] = 32'h54547280,
        RAM[1591] = 32'h25e63874,
        RAM[1592] = 32'h085574d1,
        RAM[1593] = 32'h3875900c,
        RAM[1594] = 32'h893d0d04,
        RAM[1595] = 32'h7351762d,
        RAM[1596] = 32'h75900807,
        RAM[1597] = 32'h80dc15ff,
        RAM[1598] = 32'h15555556,
        RAM[1599] = 32'hff9e3973,
        RAM[1600] = 32'h51762d75,
        RAM[1601] = 32'h90080780,
        RAM[1602] = 32'hdc15ff15,
        RAM[1603] = 32'h555556ca,
        RAM[1604] = 32'h39ea3d0d,
        RAM[1605] = 32'h688c1122,
        RAM[1606] = 32'h70812a81,
        RAM[1607] = 32'h06575856,
        RAM[1608] = 32'h7480e438,
        RAM[1609] = 32'h8e162270,
        RAM[1610] = 32'h902b7090,
        RAM[1611] = 32'h2c515558,
        RAM[1612] = 32'h807424b1,
        RAM[1613] = 32'h38983dc4,
        RAM[1614] = 32'h05537352,
        RAM[1615] = 32'h80cfc008,
        RAM[1616] = 32'h5192ac3f,
        RAM[1617] = 32'h800b9008,
        RAM[1618] = 32'h24973879,
        RAM[1619] = 32'h83e08006,
        RAM[1620] = 32'h547380c0,
        RAM[1621] = 32'h802e818f,
        RAM[1622] = 32'h38738280,
        RAM[1623] = 32'h802e8191,
        RAM[1624] = 32'h388c1622,
        RAM[1625] = 32'h57769080,
        RAM[1626] = 32'h0754738c,
        RAM[1627] = 32'h17238880,
        RAM[1628] = 32'h5280cfc0,
        RAM[1629] = 32'h0851819b,
        RAM[1630] = 32'h3f90089d,
        RAM[1631] = 32'h388c1622,
        RAM[1632] = 32'h82075473,
        RAM[1633] = 32'h8c172380,
        RAM[1634] = 32'hc3167077,
        RAM[1635] = 32'h0c90170c,
        RAM[1636] = 32'h810b9417,
        RAM[1637] = 32'h0c983d0d,
        RAM[1638] = 32'h0480cfc0,
        RAM[1639] = 32'h08aaab0b,
        RAM[1640] = 32'hbc120c54,
        RAM[1641] = 32'h8c162281,
        RAM[1642] = 32'h80075473,
        RAM[1643] = 32'h8c172390,
        RAM[1644] = 32'h08760c90,
        RAM[1645] = 32'h0890170c,
        RAM[1646] = 32'h88800b94,
        RAM[1647] = 32'h170c7480,
        RAM[1648] = 32'h2ed3388e,
        RAM[1649] = 32'h16227090,
        RAM[1650] = 32'h2b70902c,
        RAM[1651] = 32'h53555898,
        RAM[1652] = 32'ha23f9008,
        RAM[1653] = 32'h802effbd,
        RAM[1654] = 32'h388c1622,
        RAM[1655] = 32'h81075473,
        RAM[1656] = 32'h8c172398,
        RAM[1657] = 32'h3d0d0481,
        RAM[1658] = 32'h0b8c1722,
        RAM[1659] = 32'h5855fef5,
        RAM[1660] = 32'h39a81608,
        RAM[1661] = 32'h80c3922e,
        RAM[1662] = 32'h098106fe,
        RAM[1663] = 32'he4388c16,
        RAM[1664] = 32'h22888007,
        RAM[1665] = 32'h54738c17,
        RAM[1666] = 32'h2388800b,
        RAM[1667] = 32'h80cc170c,
        RAM[1668] = 32'hfedc39f3,
        RAM[1669] = 32'h3d0d7f61,
        RAM[1670] = 32'h8b1170f8,
        RAM[1671] = 32'h065c5555,
        RAM[1672] = 32'h5e729626,
        RAM[1673] = 32'h83389059,
        RAM[1674] = 32'h80792474,
        RAM[1675] = 32'h7a260753,
        RAM[1676] = 32'h80547274,
        RAM[1677] = 32'h2e098106,
        RAM[1678] = 32'h80cb387d,
        RAM[1679] = 32'h518cd93f,
        RAM[1680] = 32'h7883f726,
        RAM[1681] = 32'h80c63878,
        RAM[1682] = 32'h832a7010,
        RAM[1683] = 32'h101080d6,
        RAM[1684] = 32'hfc058c11,
        RAM[1685] = 32'h0859595a,
        RAM[1686] = 32'h76782e83,
        RAM[1687] = 32'hb0388417,
        RAM[1688] = 32'h08fc0656,
        RAM[1689] = 32'h8c170888,
        RAM[1690] = 32'h1808718c,
        RAM[1691] = 32'h120c8812,
        RAM[1692] = 32'h0c587517,
        RAM[1693] = 32'h84110881,
        RAM[1694] = 32'h0784120c,
        RAM[1695] = 32'h537d518c,
        RAM[1696] = 32'h983f8817,
        RAM[1697] = 32'h5473900c,
        RAM[1698] = 32'h8f3d0d04,
        RAM[1699] = 32'h78892a79,
        RAM[1700] = 32'h832a5b53,
        RAM[1701] = 32'h72802ebf,
        RAM[1702] = 32'h3878862a,
        RAM[1703] = 32'hb8055a84,
        RAM[1704] = 32'h7327b438,
        RAM[1705] = 32'h80db135a,
        RAM[1706] = 32'h947327ab,
        RAM[1707] = 32'h38788c2a,
        RAM[1708] = 32'h80ee055a,
        RAM[1709] = 32'h80d47327,
        RAM[1710] = 32'h9e38788f,
        RAM[1711] = 32'h2a80f705,
        RAM[1712] = 32'h5a82d473,
        RAM[1713] = 32'h27913878,
        RAM[1714] = 32'h922a80fc,
        RAM[1715] = 32'h055a8ad4,
        RAM[1716] = 32'h73278438,
        RAM[1717] = 32'h80fe5a79,
        RAM[1718] = 32'h10101080,
        RAM[1719] = 32'hd6fc058c,
        RAM[1720] = 32'h11085855,
        RAM[1721] = 32'h76752ea3,
        RAM[1722] = 32'h38841708,
        RAM[1723] = 32'hfc06707a,
        RAM[1724] = 32'h31555673,
        RAM[1725] = 32'h8f2488d5,
        RAM[1726] = 32'h38738025,
        RAM[1727] = 32'hfee6388c,
        RAM[1728] = 32'h17085776,
        RAM[1729] = 32'h752e0981,
        RAM[1730] = 32'h06df3881,
        RAM[1731] = 32'h1a5a80d7,
        RAM[1732] = 32'h8c085776,
        RAM[1733] = 32'h80d7842e,
        RAM[1734] = 32'h82c03884,
        RAM[1735] = 32'h1708fc06,
        RAM[1736] = 32'h707a3155,
        RAM[1737] = 32'h56738f24,
        RAM[1738] = 32'h81f93880,
        RAM[1739] = 32'hd7840b80,
        RAM[1740] = 32'hd7900c80,
        RAM[1741] = 32'hd7840b80,
        RAM[1742] = 32'hd78c0c73,
        RAM[1743] = 32'h8025feb2,
        RAM[1744] = 32'h3883ff76,
        RAM[1745] = 32'h2783df38,
        RAM[1746] = 32'h75892a76,
        RAM[1747] = 32'h832a5553,
        RAM[1748] = 32'h72802ebf,
        RAM[1749] = 32'h3875862a,
        RAM[1750] = 32'hb8055484,
        RAM[1751] = 32'h7327b438,
        RAM[1752] = 32'h80db1354,
        RAM[1753] = 32'h947327ab,
        RAM[1754] = 32'h38758c2a,
        RAM[1755] = 32'h80ee0554,
        RAM[1756] = 32'h80d47327,
        RAM[1757] = 32'h9e38758f,
        RAM[1758] = 32'h2a80f705,
        RAM[1759] = 32'h5482d473,
        RAM[1760] = 32'h27913875,
        RAM[1761] = 32'h922a80fc,
        RAM[1762] = 32'h05548ad4,
        RAM[1763] = 32'h73278438,
        RAM[1764] = 32'h80fe5473,
        RAM[1765] = 32'h10101080,
        RAM[1766] = 32'hd6fc0588,
        RAM[1767] = 32'h11085658,
        RAM[1768] = 32'h74782e86,
        RAM[1769] = 32'hcf388415,
        RAM[1770] = 32'h08fc0653,
        RAM[1771] = 32'h7573278d,
        RAM[1772] = 32'h38881508,
        RAM[1773] = 32'h5574782e,
        RAM[1774] = 32'h098106ea,
        RAM[1775] = 32'h388c1508,
        RAM[1776] = 32'h80d6fc0b,
        RAM[1777] = 32'h84050871,
        RAM[1778] = 32'h8c1a0c76,
        RAM[1779] = 32'h881a0c78,
        RAM[1780] = 32'h88130c78,
        RAM[1781] = 32'h8c180c5d,
        RAM[1782] = 32'h58795380,
        RAM[1783] = 32'h7a2483e6,
        RAM[1784] = 32'h3872822c,
        RAM[1785] = 32'h81712b5c,
        RAM[1786] = 32'h537a7c26,
        RAM[1787] = 32'h8198387b,
        RAM[1788] = 32'h7b065372,
        RAM[1789] = 32'h82f13879,
        RAM[1790] = 32'hfc068405,
        RAM[1791] = 32'h5a7a1070,
        RAM[1792] = 32'h7d06545b,
        RAM[1793] = 32'h7282e038,
        RAM[1794] = 32'h841a5af1,
        RAM[1795] = 32'h3988178c,
        RAM[1796] = 32'h11085858,
        RAM[1797] = 32'h76782e09,
        RAM[1798] = 32'h8106fcc2,
        RAM[1799] = 32'h38821a5a,
        RAM[1800] = 32'hfdec3978,
        RAM[1801] = 32'h17798107,
        RAM[1802] = 32'h84190c70,
        RAM[1803] = 32'h80d7900c,
        RAM[1804] = 32'h7080d78c,
        RAM[1805] = 32'h0c80d784,
        RAM[1806] = 32'h0b8c120c,
        RAM[1807] = 32'h8c110888,
        RAM[1808] = 32'h120c7481,
        RAM[1809] = 32'h0784120c,
        RAM[1810] = 32'h74117571,
        RAM[1811] = 32'h0c51537d,
        RAM[1812] = 32'h5188c63f,
        RAM[1813] = 32'h881754fc,
        RAM[1814] = 32'hac3980d6,
        RAM[1815] = 32'hfc0b8405,
        RAM[1816] = 32'h087a545c,
        RAM[1817] = 32'h798025fe,
        RAM[1818] = 32'hf83882da,
        RAM[1819] = 32'h397a097c,
        RAM[1820] = 32'h067080d6,
        RAM[1821] = 32'hfc0b8405,
        RAM[1822] = 32'h0c5c7a10,
        RAM[1823] = 32'h5b7a7c26,
        RAM[1824] = 32'h85387a85,
        RAM[1825] = 32'hb83880d6,
        RAM[1826] = 32'hfc0b8805,
        RAM[1827] = 32'h08708412,
        RAM[1828] = 32'h08fc0670,
        RAM[1829] = 32'h7c317c72,
        RAM[1830] = 32'h268f7225,
        RAM[1831] = 32'h0757575c,
        RAM[1832] = 32'h5d557280,
        RAM[1833] = 32'h2e80db38,
        RAM[1834] = 32'h797a1680,
        RAM[1835] = 32'hd6f4081b,
        RAM[1836] = 32'h90115a55,
        RAM[1837] = 32'h575b80d6,
        RAM[1838] = 32'hf008ff2e,
        RAM[1839] = 32'h8838a08f,
        RAM[1840] = 32'h13e08006,
        RAM[1841] = 32'h5776527d,
        RAM[1842] = 32'h5187cf3f,
        RAM[1843] = 32'h90085490,
        RAM[1844] = 32'h08ff2e90,
        RAM[1845] = 32'h38900876,
        RAM[1846] = 32'h27829938,
        RAM[1847] = 32'h7480d6fc,
        RAM[1848] = 32'h2e829138,
        RAM[1849] = 32'h80d6fc0b,
        RAM[1850] = 32'h88050855,
        RAM[1851] = 32'h841508fc,
        RAM[1852] = 32'h06707a31,
        RAM[1853] = 32'h7a72268f,
        RAM[1854] = 32'h72250752,
        RAM[1855] = 32'h55537283,
        RAM[1856] = 32'he6387479,
        RAM[1857] = 32'h81078417,
        RAM[1858] = 32'h0c791670,
        RAM[1859] = 32'h80d6fc0b,
        RAM[1860] = 32'h88050c75,
        RAM[1861] = 32'h81078412,
        RAM[1862] = 32'h0c547e52,
        RAM[1863] = 32'h5786fa3f,
        RAM[1864] = 32'h881754fa,
        RAM[1865] = 32'he0397583,
        RAM[1866] = 32'h2a705454,
        RAM[1867] = 32'h80742481,
        RAM[1868] = 32'h9b387282,
        RAM[1869] = 32'h2c81712b,
        RAM[1870] = 32'h80d78008,
        RAM[1871] = 32'h077080d6,
        RAM[1872] = 32'hfc0b8405,
        RAM[1873] = 32'h0c751010,
        RAM[1874] = 32'h1080d6fc,
        RAM[1875] = 32'h05881108,
        RAM[1876] = 32'h585a5d53,
        RAM[1877] = 32'h778c180c,
        RAM[1878] = 32'h7488180c,
        RAM[1879] = 32'h7688190c,
        RAM[1880] = 32'h768c160c,
        RAM[1881] = 32'hfcf33979,
        RAM[1882] = 32'h7a101010,
        RAM[1883] = 32'h80d6fc05,
        RAM[1884] = 32'h7057595d,
        RAM[1885] = 32'h8c150857,
        RAM[1886] = 32'h76752ea3,
        RAM[1887] = 32'h38841708,
        RAM[1888] = 32'hfc06707a,
        RAM[1889] = 32'h31555673,
        RAM[1890] = 32'h8f2483ca,
        RAM[1891] = 32'h38738025,
        RAM[1892] = 32'h8481388c,
        RAM[1893] = 32'h17085776,
        RAM[1894] = 32'h752e0981,
        RAM[1895] = 32'h06df3888,
        RAM[1896] = 32'h15811b70,
        RAM[1897] = 32'h8306555b,
        RAM[1898] = 32'h5572c938,
        RAM[1899] = 32'h7c830653,
        RAM[1900] = 32'h72802efd,
        RAM[1901] = 32'hb838ff1d,
        RAM[1902] = 32'hf819595d,
        RAM[1903] = 32'h88180878,
        RAM[1904] = 32'h2eea38fd,
        RAM[1905] = 32'hb539831a,
        RAM[1906] = 32'h53fc9639,
        RAM[1907] = 32'h83147082,
        RAM[1908] = 32'h2c81712b,
        RAM[1909] = 32'h80d78008,
        RAM[1910] = 32'h077080d6,
        RAM[1911] = 32'hfc0b8405,
        RAM[1912] = 32'h0c761010,
        RAM[1913] = 32'h1080d6fc,
        RAM[1914] = 32'h05881108,
        RAM[1915] = 32'h595b5e51,
        RAM[1916] = 32'h53fee139,
        RAM[1917] = 32'h80d6c008,
        RAM[1918] = 32'h17589008,
        RAM[1919] = 32'h762e818d,
        RAM[1920] = 32'h3880d6f0,
        RAM[1921] = 32'h08ff2e83,
        RAM[1922] = 32'hec387376,
        RAM[1923] = 32'h311880d6,
        RAM[1924] = 32'hc00c7387,
        RAM[1925] = 32'h06705753,
        RAM[1926] = 32'h72802e88,
        RAM[1927] = 32'h38887331,
        RAM[1928] = 32'h70155556,
        RAM[1929] = 32'h76149fff,
        RAM[1930] = 32'h06a08071,
        RAM[1931] = 32'h31177054,
        RAM[1932] = 32'h7f535753,
        RAM[1933] = 32'h84e43f90,
        RAM[1934] = 32'h08539008,
        RAM[1935] = 32'hff2e81a0,
        RAM[1936] = 32'h3880d6c0,
        RAM[1937] = 32'h08167080,
        RAM[1938] = 32'hd6c00c74,
        RAM[1939] = 32'h7580d6fc,
        RAM[1940] = 32'h0b88050c,
        RAM[1941] = 32'h74763118,
        RAM[1942] = 32'h70810751,
        RAM[1943] = 32'h5556587b,
        RAM[1944] = 32'h80d6fc2e,
        RAM[1945] = 32'h839c3879,
        RAM[1946] = 32'h8f2682cb,
        RAM[1947] = 32'h38810b84,
        RAM[1948] = 32'h150c8415,
        RAM[1949] = 32'h08fc0670,
        RAM[1950] = 32'h7a317a72,
        RAM[1951] = 32'h268f7225,
        RAM[1952] = 32'h07525553,
        RAM[1953] = 32'h72802efc,
        RAM[1954] = 32'hf93880db,
        RAM[1955] = 32'h3990089f,
        RAM[1956] = 32'hff065372,
        RAM[1957] = 32'hfeeb3877,
        RAM[1958] = 32'h80d6c00c,
        RAM[1959] = 32'h80d6fc0b,
        RAM[1960] = 32'h8805087b,
        RAM[1961] = 32'h18810784,
        RAM[1962] = 32'h120c5580,
        RAM[1963] = 32'hd6ec0878,
        RAM[1964] = 32'h27863877,
        RAM[1965] = 32'h80d6ec0c,
        RAM[1966] = 32'h80d6e808,
        RAM[1967] = 32'h7827fcac,
        RAM[1968] = 32'h387780d6,
        RAM[1969] = 32'he80c8415,
        RAM[1970] = 32'h08fc0670,
        RAM[1971] = 32'h7a317a72,
        RAM[1972] = 32'h268f7225,
        RAM[1973] = 32'h07525553,
        RAM[1974] = 32'h72802efc,
        RAM[1975] = 32'ha5388839,
        RAM[1976] = 32'h80745456,
        RAM[1977] = 32'hfedb397d,
        RAM[1978] = 32'h5183ae3f,
        RAM[1979] = 32'h800b900c,
        RAM[1980] = 32'h8f3d0d04,
        RAM[1981] = 32'h73538074,
        RAM[1982] = 32'h24a93872,
        RAM[1983] = 32'h822c8171,
        RAM[1984] = 32'h2b80d780,
        RAM[1985] = 32'h08077080,
        RAM[1986] = 32'hd6fc0b84,
        RAM[1987] = 32'h050c5d53,
        RAM[1988] = 32'h778c180c,
        RAM[1989] = 32'h7488180c,
        RAM[1990] = 32'h7688190c,
        RAM[1991] = 32'h768c160c,
        RAM[1992] = 32'hf9b73983,
        RAM[1993] = 32'h1470822c,
        RAM[1994] = 32'h81712b80,
        RAM[1995] = 32'hd7800807,
        RAM[1996] = 32'h7080d6fc,
        RAM[1997] = 32'h0b84050c,
        RAM[1998] = 32'h5e5153d4,
        RAM[1999] = 32'h397b7b06,
        RAM[2000] = 32'h5372fca3,
        RAM[2001] = 32'h38841a7b,
        RAM[2002] = 32'h105c5af1,
        RAM[2003] = 32'h39ff1a81,
        RAM[2004] = 32'h11515af7,
        RAM[2005] = 32'hb9397817,
        RAM[2006] = 32'h79810784,
        RAM[2007] = 32'h190c8c18,
        RAM[2008] = 32'h08881908,
        RAM[2009] = 32'h718c120c,
        RAM[2010] = 32'h88120c59,
        RAM[2011] = 32'h7080d790,
        RAM[2012] = 32'h0c7080d7,
        RAM[2013] = 32'h8c0c80d7,
        RAM[2014] = 32'h840b8c12,
        RAM[2015] = 32'h0c8c1108,
        RAM[2016] = 32'h88120c74,
        RAM[2017] = 32'h81078412,
        RAM[2018] = 32'h0c741175,
        RAM[2019] = 32'h710c5153,
        RAM[2020] = 32'hf9bd3975,
        RAM[2021] = 32'h17841108,
        RAM[2022] = 32'h81078412,
        RAM[2023] = 32'h0c538c17,
        RAM[2024] = 32'h08881808,
        RAM[2025] = 32'h718c120c,
        RAM[2026] = 32'h88120c58,
        RAM[2027] = 32'h7d5181e9,
        RAM[2028] = 32'h3f881754,
        RAM[2029] = 32'hf5cf3972,
        RAM[2030] = 32'h84150cf4,
        RAM[2031] = 32'h1af80670,
        RAM[2032] = 32'h841e0881,
        RAM[2033] = 32'h0607841e,
        RAM[2034] = 32'h0c701d54,
        RAM[2035] = 32'h5b850b84,
        RAM[2036] = 32'h140c850b,
        RAM[2037] = 32'h88140c8f,
        RAM[2038] = 32'h7b27fdcf,
        RAM[2039] = 32'h38881c52,
        RAM[2040] = 32'h7d51ec9e,
        RAM[2041] = 32'h3f80d6fc,
        RAM[2042] = 32'h0b880508,
        RAM[2043] = 32'h80d6c008,
        RAM[2044] = 32'h5955fdb7,
        RAM[2045] = 32'h397780d6,
        RAM[2046] = 32'hc00c7380,
        RAM[2047] = 32'hd6f00cfc,
        RAM[2048] = 32'h91397284,
        RAM[2049] = 32'h150cfda3,
        RAM[2050] = 32'h39fc3d0d,
        RAM[2051] = 32'h76797102,
        RAM[2052] = 32'h8c059f05,
        RAM[2053] = 32'h33575553,
        RAM[2054] = 32'h55837227,
        RAM[2055] = 32'h8a387483,
        RAM[2056] = 32'h06517080,
        RAM[2057] = 32'h2ea238ff,
        RAM[2058] = 32'h125271ff,
        RAM[2059] = 32'h2e933873,
        RAM[2060] = 32'h73708105,
        RAM[2061] = 32'h5534ff12,
        RAM[2062] = 32'h5271ff2e,
        RAM[2063] = 32'h098106ef,
        RAM[2064] = 32'h3874900c,
        RAM[2065] = 32'h863d0d04,
        RAM[2066] = 32'h7474882b,
        RAM[2067] = 32'h75077071,
        RAM[2068] = 32'h902b0751,
        RAM[2069] = 32'h54518f72,
        RAM[2070] = 32'h27a53872,
        RAM[2071] = 32'h71708405,
        RAM[2072] = 32'h530c7271,
        RAM[2073] = 32'h70840553,
        RAM[2074] = 32'h0c727170,
        RAM[2075] = 32'h8405530c,
        RAM[2076] = 32'h72717084,
        RAM[2077] = 32'h05530cf0,
        RAM[2078] = 32'h1252718f,
        RAM[2079] = 32'h26dd3883,
        RAM[2080] = 32'h72279038,
        RAM[2081] = 32'h72717084,
        RAM[2082] = 32'h05530cfc,
        RAM[2083] = 32'h12527183,
        RAM[2084] = 32'h26f23870,
        RAM[2085] = 32'h53ff9039,
        RAM[2086] = 32'h0404fd3d,
        RAM[2087] = 32'h0d800b80,
        RAM[2088] = 32'hdfb40c76,
        RAM[2089] = 32'h5184ee3f,
        RAM[2090] = 32'h90085390,
        RAM[2091] = 32'h08ff2e88,
        RAM[2092] = 32'h3872900c,
        RAM[2093] = 32'h853d0d04,
        RAM[2094] = 32'h80dfb408,
        RAM[2095] = 32'h5473802e,
        RAM[2096] = 32'hf0387574,
        RAM[2097] = 32'h710c5272,
        RAM[2098] = 32'h900c853d,
        RAM[2099] = 32'h0d04f93d,
        RAM[2100] = 32'h0d797c55,
        RAM[2101] = 32'h7b548e11,
        RAM[2102] = 32'h2270902b,
        RAM[2103] = 32'h70902c55,
        RAM[2104] = 32'h5780cfc0,
        RAM[2105] = 32'h08535856,
        RAM[2106] = 32'h83f33f90,
        RAM[2107] = 32'h0857800b,
        RAM[2108] = 32'h90082493,
        RAM[2109] = 32'h3880d016,
        RAM[2110] = 32'h08900805,
        RAM[2111] = 32'h80d0170c,
        RAM[2112] = 32'h76900c89,
        RAM[2113] = 32'h3d0d048c,
        RAM[2114] = 32'h162283df,
        RAM[2115] = 32'hff065574,
        RAM[2116] = 32'h8c172376,
        RAM[2117] = 32'h900c893d,
        RAM[2118] = 32'h0d04fa3d,
        RAM[2119] = 32'h0d788c11,
        RAM[2120] = 32'h2270882a,
        RAM[2121] = 32'h70810651,
        RAM[2122] = 32'h57585674,
        RAM[2123] = 32'ha9388c16,
        RAM[2124] = 32'h2283dfff,
        RAM[2125] = 32'h0655748c,
        RAM[2126] = 32'h17237a54,
        RAM[2127] = 32'h79538e16,
        RAM[2128] = 32'h2270902b,
        RAM[2129] = 32'h70902c54,
        RAM[2130] = 32'h5680cfc0,
        RAM[2131] = 32'h08525681,
        RAM[2132] = 32'hb23f883d,
        RAM[2133] = 32'h0d048254,
        RAM[2134] = 32'h80538e16,
        RAM[2135] = 32'h2270902b,
        RAM[2136] = 32'h70902c54,
        RAM[2137] = 32'h5680cfc0,
        RAM[2138] = 32'h08525782,
        RAM[2139] = 32'hb83f8c16,
        RAM[2140] = 32'h2283dfff,
        RAM[2141] = 32'h0655748c,
        RAM[2142] = 32'h17237a54,
        RAM[2143] = 32'h79538e16,
        RAM[2144] = 32'h2270902b,
        RAM[2145] = 32'h70902c54,
        RAM[2146] = 32'h5680cfc0,
        RAM[2147] = 32'h08525680,
        RAM[2148] = 32'hf23f883d,
        RAM[2149] = 32'h0d04f93d,
        RAM[2150] = 32'h0d797c55,
        RAM[2151] = 32'h7b548e11,
        RAM[2152] = 32'h2270902b,
        RAM[2153] = 32'h70902c55,
        RAM[2154] = 32'h5780cfc0,
        RAM[2155] = 32'h08535856,
        RAM[2156] = 32'h81f33f90,
        RAM[2157] = 32'h08579008,
        RAM[2158] = 32'hff2e9938,
        RAM[2159] = 32'h8c1622a0,
        RAM[2160] = 32'h80075574,
        RAM[2161] = 32'h8c172390,
        RAM[2162] = 32'h0880d017,
        RAM[2163] = 32'h0c76900c,
        RAM[2164] = 32'h893d0d04,
        RAM[2165] = 32'h8c162283,
        RAM[2166] = 32'hdfff0655,
        RAM[2167] = 32'h748c1723,
        RAM[2168] = 32'h76900c89,
        RAM[2169] = 32'h3d0d04fe,
        RAM[2170] = 32'h3d0d748e,
        RAM[2171] = 32'h11227090,
        RAM[2172] = 32'h2b70902c,
        RAM[2173] = 32'h55515153,
        RAM[2174] = 32'h80cfc008,
        RAM[2175] = 32'h51bd3f84,
        RAM[2176] = 32'h3d0d04fb,
        RAM[2177] = 32'h3d0d800b,
        RAM[2178] = 32'h80dfb40c,
        RAM[2179] = 32'h7a537952,
        RAM[2180] = 32'h785182f9,
        RAM[2181] = 32'h3f900855,
        RAM[2182] = 32'h9008ff2e,
        RAM[2183] = 32'h88387490,
        RAM[2184] = 32'h0c873d0d,
        RAM[2185] = 32'h0480dfb4,
        RAM[2186] = 32'h08567580,
        RAM[2187] = 32'h2ef03877,
        RAM[2188] = 32'h76710c54,
        RAM[2189] = 32'h74900c87,
        RAM[2190] = 32'h3d0d04fd,
        RAM[2191] = 32'h3d0d800b,
        RAM[2192] = 32'h80dfb40c,
        RAM[2193] = 32'h765184c4,
        RAM[2194] = 32'h3f900853,
        RAM[2195] = 32'h9008ff2e,
        RAM[2196] = 32'h88387290,
        RAM[2197] = 32'h0c853d0d,
        RAM[2198] = 32'h0480dfb4,
        RAM[2199] = 32'h08547380,
        RAM[2200] = 32'h2ef03875,
        RAM[2201] = 32'h74710c52,
        RAM[2202] = 32'h72900c85,
        RAM[2203] = 32'h3d0d04fc,
        RAM[2204] = 32'h3d0d800b,
        RAM[2205] = 32'h80dfb40c,
        RAM[2206] = 32'h78527751,
        RAM[2207] = 32'h86ac3f90,
        RAM[2208] = 32'h08549008,
        RAM[2209] = 32'hff2e8838,
        RAM[2210] = 32'h73900c86,
        RAM[2211] = 32'h3d0d0480,
        RAM[2212] = 32'hdfb40855,
        RAM[2213] = 32'h74802ef0,
        RAM[2214] = 32'h38767571,
        RAM[2215] = 32'h0c537390,
        RAM[2216] = 32'h0c863d0d,
        RAM[2217] = 32'h04fb3d0d,
        RAM[2218] = 32'h800b80df,
        RAM[2219] = 32'hb40c7a53,
        RAM[2220] = 32'h79527851,
        RAM[2221] = 32'h84883f90,
        RAM[2222] = 32'h08559008,
        RAM[2223] = 32'hff2e8838,
        RAM[2224] = 32'h74900c87,
        RAM[2225] = 32'h3d0d0480,
        RAM[2226] = 32'hdfb40856,
        RAM[2227] = 32'h75802ef0,
        RAM[2228] = 32'h38777671,
        RAM[2229] = 32'h0c547490,
        RAM[2230] = 32'h0c873d0d,
        RAM[2231] = 32'h04fb3d0d,
        RAM[2232] = 32'h800b80df,
        RAM[2233] = 32'hb40c7a53,
        RAM[2234] = 32'h79527851,
        RAM[2235] = 32'h82933f90,
        RAM[2236] = 32'h08559008,
        RAM[2237] = 32'hff2e8838,
        RAM[2238] = 32'h74900c87,
        RAM[2239] = 32'h3d0d0480,
        RAM[2240] = 32'hdfb40856,
        RAM[2241] = 32'h75802ef0,
        RAM[2242] = 32'h38777671,
        RAM[2243] = 32'h0c547490,
        RAM[2244] = 32'h0c873d0d,
        RAM[2245] = 32'h04fe3d0d,
        RAM[2246] = 32'h80dfac08,
        RAM[2247] = 32'h51708a38,
        RAM[2248] = 32'h80dfb870,
        RAM[2249] = 32'h80dfac0c,
        RAM[2250] = 32'h51707512,
        RAM[2251] = 32'h5252ff53,
        RAM[2252] = 32'h7087fb80,
        RAM[2253] = 32'h80268838,
        RAM[2254] = 32'h7080dfac,
        RAM[2255] = 32'h0c715372,
        RAM[2256] = 32'h900c843d,
        RAM[2257] = 32'h0d04fd3d,
        RAM[2258] = 32'h0d800b80,
        RAM[2259] = 32'hceb40854,
        RAM[2260] = 32'h5472812e,
        RAM[2261] = 32'h9b387380,
        RAM[2262] = 32'hdfb00cc2,
        RAM[2263] = 32'hfd3fc1a4,
        RAM[2264] = 32'h3f80df84,
        RAM[2265] = 32'h528151c5,
        RAM[2266] = 32'h9e3f9008,
        RAM[2267] = 32'h5185bb3f,
        RAM[2268] = 32'h7280dfb0,
        RAM[2269] = 32'h0cc2e33f,
        RAM[2270] = 32'hc18a3f80,
        RAM[2271] = 32'hdf845281,
        RAM[2272] = 32'h51c5843f,
        RAM[2273] = 32'h90085185,
        RAM[2274] = 32'ha13f00ff,
        RAM[2275] = 32'h39f53d0d,
        RAM[2276] = 32'h7e6080df,
        RAM[2277] = 32'hb008705b,
        RAM[2278] = 32'h585b5b75,
        RAM[2279] = 32'h80c23877,
        RAM[2280] = 32'h7a25a138,
        RAM[2281] = 32'h771b7033,
        RAM[2282] = 32'h7081ff06,
        RAM[2283] = 32'h58585975,
        RAM[2284] = 32'h8a2e9838,
        RAM[2285] = 32'h7681ff06,
        RAM[2286] = 32'h51c1fe3f,
        RAM[2287] = 32'h81185879,
        RAM[2288] = 32'h7824e138,
        RAM[2289] = 32'h79900c8d,
        RAM[2290] = 32'h3d0d048d,
        RAM[2291] = 32'h51c1ea3f,
        RAM[2292] = 32'h78337081,
        RAM[2293] = 32'hff065257,
        RAM[2294] = 32'hc1df3f81,
        RAM[2295] = 32'h1858e039,
        RAM[2296] = 32'h79557a54,
        RAM[2297] = 32'h7d538552,
        RAM[2298] = 32'h8d3dfc05,
        RAM[2299] = 32'h51c0d73f,
        RAM[2300] = 32'h90085684,
        RAM[2301] = 32'hae3f7b90,
        RAM[2302] = 32'h080c7590,
        RAM[2303] = 32'h0c8d3d0d,
        RAM[2304] = 32'h04f63d0d,
        RAM[2305] = 32'h7d7f80df,
        RAM[2306] = 32'hb008705b,
        RAM[2307] = 32'h585a5a75,
        RAM[2308] = 32'h80c13877,
        RAM[2309] = 32'h7925b338,
        RAM[2310] = 32'hc0fa3f90,
        RAM[2311] = 32'h0881ff06,
        RAM[2312] = 32'h708d3270,
        RAM[2313] = 32'h30709f2a,
        RAM[2314] = 32'h51515757,
        RAM[2315] = 32'h768a2e80,
        RAM[2316] = 32'hc4387580,
        RAM[2317] = 32'h2ebf3877,
        RAM[2318] = 32'h1a567676,
        RAM[2319] = 32'h347651c0,
        RAM[2320] = 32'hf83f8118,
        RAM[2321] = 32'h58787824,
        RAM[2322] = 32'hcf387756,
        RAM[2323] = 32'h75900c8c,
        RAM[2324] = 32'h3d0d0478,
        RAM[2325] = 32'h5579547c,
        RAM[2326] = 32'h5384528c,
        RAM[2327] = 32'h3dfc0551,
        RAM[2328] = 32'hffbfe33f,
        RAM[2329] = 32'h90085683,
        RAM[2330] = 32'hba3f7a90,
        RAM[2331] = 32'h080c7590,
        RAM[2332] = 32'h0c8c3d0d,
        RAM[2333] = 32'h04771a56,
        RAM[2334] = 32'h8a763481,
        RAM[2335] = 32'h18588d51,
        RAM[2336] = 32'hc0b73f8a,
        RAM[2337] = 32'h51c0b23f,
        RAM[2338] = 32'h7756c139,
        RAM[2339] = 32'hfb3d0d80,
        RAM[2340] = 32'hdfb00870,
        RAM[2341] = 32'h56547388,
        RAM[2342] = 32'h3874900c,
        RAM[2343] = 32'h873d0d04,
        RAM[2344] = 32'h77538352,
        RAM[2345] = 32'h873dfc05,
        RAM[2346] = 32'h51ffbf9a,
        RAM[2347] = 32'h3f900854,
        RAM[2348] = 32'h82f13f75,
        RAM[2349] = 32'h90080c73,
        RAM[2350] = 32'h900c873d,
        RAM[2351] = 32'h0d04fa3d,
        RAM[2352] = 32'h0d80dfb0,
        RAM[2353] = 32'h08802ea3,
        RAM[2354] = 32'h387a5579,
        RAM[2355] = 32'h54785386,
        RAM[2356] = 32'h52883dfc,
        RAM[2357] = 32'h0551ffbe,
        RAM[2358] = 32'hed3f9008,
        RAM[2359] = 32'h5682c43f,
        RAM[2360] = 32'h7690080c,
        RAM[2361] = 32'h75900c88,
        RAM[2362] = 32'h3d0d0482,
        RAM[2363] = 32'hb63f9d0b,
        RAM[2364] = 32'h90080cff,
        RAM[2365] = 32'h0b900c88,
        RAM[2366] = 32'h3d0d04fb,
        RAM[2367] = 32'h3d0d7779,
        RAM[2368] = 32'h56568070,
        RAM[2369] = 32'h54547375,
        RAM[2370] = 32'h259f3874,
        RAM[2371] = 32'h101010f8,
        RAM[2372] = 32'h05527216,
        RAM[2373] = 32'h70337074,
        RAM[2374] = 32'h2b760781,
        RAM[2375] = 32'h16f81656,
        RAM[2376] = 32'h56565151,
        RAM[2377] = 32'h747324ea,
        RAM[2378] = 32'h3873900c,
        RAM[2379] = 32'h873d0d04,
        RAM[2380] = 32'hfc3d0d76,
        RAM[2381] = 32'h785555bc,
        RAM[2382] = 32'h53805273,
        RAM[2383] = 32'h51f5ca3f,
        RAM[2384] = 32'h84527451,
        RAM[2385] = 32'hffb53f90,
        RAM[2386] = 32'h08742384,
        RAM[2387] = 32'h52841551,
        RAM[2388] = 32'hffa93f90,
        RAM[2389] = 32'h08821523,
        RAM[2390] = 32'h84528815,
        RAM[2391] = 32'h51ff9c3f,
        RAM[2392] = 32'h90088415,
        RAM[2393] = 32'h0c84528c,
        RAM[2394] = 32'h1551ff8f,
        RAM[2395] = 32'h3f900888,
        RAM[2396] = 32'h15238452,
        RAM[2397] = 32'h901551ff,
        RAM[2398] = 32'h823f9008,
        RAM[2399] = 32'h8a152384,
        RAM[2400] = 32'h52941551,
        RAM[2401] = 32'hfef53f90,
        RAM[2402] = 32'h088c1523,
        RAM[2403] = 32'h84529815,
        RAM[2404] = 32'h51fee83f,
        RAM[2405] = 32'h90088e15,
        RAM[2406] = 32'h2388529c,
        RAM[2407] = 32'h1551fedb,
        RAM[2408] = 32'h3f900890,
        RAM[2409] = 32'h150c863d,
        RAM[2410] = 32'h0d04e93d,
        RAM[2411] = 32'h0d6a80df,
        RAM[2412] = 32'hb0085757,
        RAM[2413] = 32'h75933880,
        RAM[2414] = 32'hc0800b84,
        RAM[2415] = 32'h180c75ac,
        RAM[2416] = 32'h180c7590,
        RAM[2417] = 32'h0c993d0d,
        RAM[2418] = 32'h04893d70,
        RAM[2419] = 32'h556a5455,
        RAM[2420] = 32'h8a52993d,
        RAM[2421] = 32'hffbc0551,
        RAM[2422] = 32'hffbceb3f,
        RAM[2423] = 32'h90087753,
        RAM[2424] = 32'h755256fe,
        RAM[2425] = 32'hcb3fbc3f,
        RAM[2426] = 32'h7790080c,
        RAM[2427] = 32'h75900c99,
        RAM[2428] = 32'h3d0d04fc,
        RAM[2429] = 32'h3d0d8154,
        RAM[2430] = 32'h80dfb008,
        RAM[2431] = 32'h88387390,
        RAM[2432] = 32'h0c863d0d,
        RAM[2433] = 32'h04765397,
        RAM[2434] = 32'hb952863d,
        RAM[2435] = 32'hfc0551ff,
        RAM[2436] = 32'hbcb43f90,
        RAM[2437] = 32'h08548c3f,
        RAM[2438] = 32'h7490080c,
        RAM[2439] = 32'h73900c86,
        RAM[2440] = 32'h3d0d0480,
        RAM[2441] = 32'hcfc00890,
        RAM[2442] = 32'h0c04f73d,
        RAM[2443] = 32'h0d7b80cf,
        RAM[2444] = 32'hc00882c8,
        RAM[2445] = 32'h11085a54,
        RAM[2446] = 32'h5a77802e,
        RAM[2447] = 32'h80da3881,
        RAM[2448] = 32'h88188419,
        RAM[2449] = 32'h08ff0581,
        RAM[2450] = 32'h712b5955,
        RAM[2451] = 32'h59807424,
        RAM[2452] = 32'h80ea3880,
        RAM[2453] = 32'h7424b538,
        RAM[2454] = 32'h73822b78,
        RAM[2455] = 32'h11880556,
        RAM[2456] = 32'h56818019,
        RAM[2457] = 32'h08770653,
        RAM[2458] = 32'h72802eb6,
        RAM[2459] = 32'h38781670,
        RAM[2460] = 32'h08535379,
        RAM[2461] = 32'h51740853,
        RAM[2462] = 32'h722dff14,
        RAM[2463] = 32'hfc17fc17,
        RAM[2464] = 32'h79812c5a,
        RAM[2465] = 32'h57575473,
        RAM[2466] = 32'h8025d638,
        RAM[2467] = 32'h77085877,
        RAM[2468] = 32'hffad3880,
        RAM[2469] = 32'hcfc00853,
        RAM[2470] = 32'hbc1308a5,
        RAM[2471] = 32'h387951f9,
        RAM[2472] = 32'he93f7408,
        RAM[2473] = 32'h53722dff,
        RAM[2474] = 32'h14fc17fc,
        RAM[2475] = 32'h1779812c,
        RAM[2476] = 32'h5a575754,
        RAM[2477] = 32'h738025ff,
        RAM[2478] = 32'ha838d139,
        RAM[2479] = 32'h8057ff93,
        RAM[2480] = 32'h397251bc,
        RAM[2481] = 32'h13085372,
        RAM[2482] = 32'h2d7951f9,
        RAM[2483] = 32'hbd3fff3d,
        RAM[2484] = 32'h0d80df8c,
        RAM[2485] = 32'h0bfc0570,
        RAM[2486] = 32'h08525270,
        RAM[2487] = 32'hff2e9138,
        RAM[2488] = 32'h702dfc12,
        RAM[2489] = 32'h70085252,
        RAM[2490] = 32'h70ff2e09,
        RAM[2491] = 32'h8106f138,
        RAM[2492] = 32'h833d0d04,
        RAM[2493] = 32'h04ffbccd,
        RAM[2494] = 32'h3f040000,
        RAM[2495] = 32'h00ffffff,
        RAM[2496] = 32'hff00ffff,
        RAM[2497] = 32'hffff00ff,
        RAM[2498] = 32'hffffff00,
        RAM[2499] = 32'h00000064,
        RAM[2500] = 32'h0a696e74,
        RAM[2501] = 32'h65727275,
        RAM[2502] = 32'h70742074,
        RAM[2503] = 32'h696d6572,
        RAM[2504] = 32'h0a000000,
        RAM[2505] = 32'h43000000,
        RAM[2506] = 32'h64756d6d,
        RAM[2507] = 32'h792e6578,
        RAM[2508] = 32'h65000000,
        RAM[2509] = 32'h00000000,
        RAM[2510] = 32'h00000000,
        RAM[2511] = 32'h00000000,
        RAM[2512] = 32'h00002f94,
        RAM[2513] = 32'h000005b9,
        RAM[2514] = 32'h000005cf,
        RAM[2515] = 32'h000005a6,
        RAM[2516] = 32'h000005b0,
        RAM[2517] = 32'h000005a6,
        RAM[2518] = 32'h000005a6,
        RAM[2519] = 32'h000005a6,
        RAM[2520] = 32'h000005a6,
        RAM[2521] = 32'h000005a6,
        RAM[2522] = 32'h000005a6,
        RAM[2523] = 32'h000005a6,
        RAM[2524] = 32'h000005a6,
        RAM[2525] = 32'h000005a6,
        RAM[2526] = 32'h000005a6,
        RAM[2527] = 32'h000005a6,
        RAM[2528] = 32'h000005a6,
        RAM[2529] = 32'h000005a6,
        RAM[2530] = 32'h000005a6,
        RAM[2531] = 32'h000005a6,
        RAM[2532] = 32'h000005a6,
        RAM[2533] = 32'h000005a6,
        RAM[2534] = 32'h000005a6,
        RAM[2535] = 32'h000005a6,
        RAM[2536] = 32'h000005a6,
        RAM[2537] = 32'h000005a6,
        RAM[2538] = 32'h000005a6,
        RAM[2539] = 32'h000005a6,
        RAM[2540] = 32'h000005a6,
        RAM[2541] = 32'h000005a6,
        RAM[2542] = 32'h000005a6,
        RAM[2543] = 32'h000005a6,
        RAM[2544] = 32'h000005a6,
        RAM[2545] = 32'h000027c4,
        RAM[2546] = 32'h00000000,
        RAM[2547] = 32'h00002a2c,
        RAM[2548] = 32'h00002a88,
        RAM[2549] = 32'h00002ae4,
        RAM[2550] = 32'h00000000,
        RAM[2551] = 32'h00000000,
        RAM[2552] = 32'h00000000,
        RAM[2553] = 32'h00000000,
        RAM[2554] = 32'h00000000,
        RAM[2555] = 32'h00000000,
        RAM[2556] = 32'h00000000,
        RAM[2557] = 32'h00000000,
        RAM[2558] = 32'h00000000,
        RAM[2559] = 32'h00002720,
        RAM[2560] = 32'h00000000,
        RAM[2561] = 32'h00000000,
        RAM[2562] = 32'h00000000,
        RAM[2563] = 32'h00000000,
        RAM[2564] = 32'h00000000,
        RAM[2565] = 32'h00000000,
        RAM[2566] = 32'h00000000,
        RAM[2567] = 32'h00000000,
        RAM[2568] = 32'h00000000,
        RAM[2569] = 32'h00000000,
        RAM[2570] = 32'h00000000,
        RAM[2571] = 32'h00000000,
        RAM[2572] = 32'h00000000,
        RAM[2573] = 32'h00000000,
        RAM[2574] = 32'h00000000,
        RAM[2575] = 32'h00000000,
        RAM[2576] = 32'h00000000,
        RAM[2577] = 32'h00000000,
        RAM[2578] = 32'h00000000,
        RAM[2579] = 32'h00000000,
        RAM[2580] = 32'h00000000,
        RAM[2581] = 32'h00000000,
        RAM[2582] = 32'h00000000,
        RAM[2583] = 32'h00000000,
        RAM[2584] = 32'h00000000,
        RAM[2585] = 32'h00000000,
        RAM[2586] = 32'h00000000,
        RAM[2587] = 32'h00000000,
        RAM[2588] = 32'h00000001,
        RAM[2589] = 32'h330eabcd,
        RAM[2590] = 32'h1234e66d,
        RAM[2591] = 32'hdeec0005,
        RAM[2592] = 32'h000b0000,
        RAM[2593] = 32'h00000000,
        RAM[2594] = 32'h00000000,
        RAM[2595] = 32'h00000000,
        RAM[2596] = 32'h00000000,
        RAM[2597] = 32'h00000000,
        RAM[2598] = 32'h00000000,
        RAM[2599] = 32'h00000000,
        RAM[2600] = 32'h00000000,
        RAM[2601] = 32'h00000000,
        RAM[2602] = 32'h00000000,
        RAM[2603] = 32'h00000000,
        RAM[2604] = 32'h00000000,
        RAM[2605] = 32'h00000000,
        RAM[2606] = 32'h00000000,
        RAM[2607] = 32'h00000000,
        RAM[2608] = 32'h00000000,
        RAM[2609] = 32'h00000000,
        RAM[2610] = 32'h00000000,
        RAM[2611] = 32'h00000000,
        RAM[2612] = 32'h00000000,
        RAM[2613] = 32'h00000000,
        RAM[2614] = 32'h00000000,
        RAM[2615] = 32'h00000000,
        RAM[2616] = 32'h00000000,
        RAM[2617] = 32'h00000000,
        RAM[2618] = 32'h00000000,
        RAM[2619] = 32'h00000000,
        RAM[2620] = 32'h00000000,
        RAM[2621] = 32'h00000000,
        RAM[2622] = 32'h00000000,
        RAM[2623] = 32'h00000000,
        RAM[2624] = 32'h00000000,
        RAM[2625] = 32'h00000000,
        RAM[2626] = 32'h00000000,
        RAM[2627] = 32'h00000000,
        RAM[2628] = 32'h00000000,
        RAM[2629] = 32'h00000000,
        RAM[2630] = 32'h00000000,
        RAM[2631] = 32'h00000000,
        RAM[2632] = 32'h00000000,
        RAM[2633] = 32'h00000000,
        RAM[2634] = 32'h00000000,
        RAM[2635] = 32'h00000000,
        RAM[2636] = 32'h00000000,
        RAM[2637] = 32'h00000000,
        RAM[2638] = 32'h00000000,
        RAM[2639] = 32'h00000000,
        RAM[2640] = 32'h00000000,
        RAM[2641] = 32'h00000000,
        RAM[2642] = 32'h00000000,
        RAM[2643] = 32'h00000000,
        RAM[2644] = 32'h00000000,
        RAM[2645] = 32'h00000000,
        RAM[2646] = 32'h00000000,
        RAM[2647] = 32'h00000000,
        RAM[2648] = 32'h00000000,
        RAM[2649] = 32'h00000000,
        RAM[2650] = 32'h00000000,
        RAM[2651] = 32'h00000000,
        RAM[2652] = 32'h00000000,
        RAM[2653] = 32'h00000000,
        RAM[2654] = 32'h00000000,
        RAM[2655] = 32'h00000000,
        RAM[2656] = 32'h00000000,
        RAM[2657] = 32'h00000000,
        RAM[2658] = 32'h00000000,
        RAM[2659] = 32'h00000000,
        RAM[2660] = 32'h00000000,
        RAM[2661] = 32'h00000000,
        RAM[2662] = 32'h00000000,
        RAM[2663] = 32'h00000000,
        RAM[2664] = 32'h00000000,
        RAM[2665] = 32'h00000000,
        RAM[2666] = 32'h00000000,
        RAM[2667] = 32'h00000000,
        RAM[2668] = 32'h00000000,
        RAM[2669] = 32'h00000000,
        RAM[2670] = 32'h00000000,
        RAM[2671] = 32'h00000000,
        RAM[2672] = 32'h00000000,
        RAM[2673] = 32'h00000000,
        RAM[2674] = 32'h00000000,
        RAM[2675] = 32'h00000000,
        RAM[2676] = 32'h00000000,
        RAM[2677] = 32'h00000000,
        RAM[2678] = 32'h00000000,
        RAM[2679] = 32'h00000000,
        RAM[2680] = 32'h00000000,
        RAM[2681] = 32'h00000000,
        RAM[2682] = 32'h00000000,
        RAM[2683] = 32'h00000000,
        RAM[2684] = 32'h00000000,
        RAM[2685] = 32'h00000000,
        RAM[2686] = 32'h00000000,
        RAM[2687] = 32'h00000000,
        RAM[2688] = 32'h00000000,
        RAM[2689] = 32'h00000000,
        RAM[2690] = 32'h00000000,
        RAM[2691] = 32'h00000000,
        RAM[2692] = 32'h00000000,
        RAM[2693] = 32'h00000000,
        RAM[2694] = 32'h00000000,
        RAM[2695] = 32'h00000000,
        RAM[2696] = 32'h00000000,
        RAM[2697] = 32'h00000000,
        RAM[2698] = 32'h00000000,
        RAM[2699] = 32'h00000000,
        RAM[2700] = 32'h00000000,
        RAM[2701] = 32'h00000000,
        RAM[2702] = 32'h00000000,
        RAM[2703] = 32'h00000000,
        RAM[2704] = 32'h00000000,
        RAM[2705] = 32'h00000000,
        RAM[2706] = 32'h00000000,
        RAM[2707] = 32'h00000000,
        RAM[2708] = 32'h00000000,
        RAM[2709] = 32'h00000000,
        RAM[2710] = 32'h00000000,
        RAM[2711] = 32'h00000000,
        RAM[2712] = 32'h00000000,
        RAM[2713] = 32'h00000000,
        RAM[2714] = 32'h00000000,
        RAM[2715] = 32'h00000000,
        RAM[2716] = 32'h00000000,
        RAM[2717] = 32'h00000000,
        RAM[2718] = 32'h00000000,
        RAM[2719] = 32'h00000000,
        RAM[2720] = 32'h00000000,
        RAM[2721] = 32'h00000000,
        RAM[2722] = 32'h00000000,
        RAM[2723] = 32'h00000000,
        RAM[2724] = 32'h00000000,
        RAM[2725] = 32'h00000000,
        RAM[2726] = 32'h00000000,
        RAM[2727] = 32'h00000000,
        RAM[2728] = 32'h00000000,
        RAM[2729] = 32'h00000000,
        RAM[2730] = 32'h00000000,
        RAM[2731] = 32'h00000000,
        RAM[2732] = 32'h00000000,
        RAM[2733] = 32'h00000000,
        RAM[2734] = 32'h00000000,
        RAM[2735] = 32'h00000000,
        RAM[2736] = 32'h00000000,
        RAM[2737] = 32'h00000000,
        RAM[2738] = 32'h00000000,
        RAM[2739] = 32'h00000000,
        RAM[2740] = 32'h00000000,
        RAM[2741] = 32'h00000000,
        RAM[2742] = 32'h00000000,
        RAM[2743] = 32'h00000000,
        RAM[2744] = 32'h00000000,
        RAM[2745] = 32'h00000000,
        RAM[2746] = 32'h00000000,
        RAM[2747] = 32'h00000000,
        RAM[2748] = 32'h00000000,
        RAM[2749] = 32'h00000000,
        RAM[2750] = 32'h00000000,
        RAM[2751] = 32'h00000000,
        RAM[2752] = 32'h00000000,
        RAM[2753] = 32'h00000000,
        RAM[2754] = 32'h00000000,
        RAM[2755] = 32'h00000000,
        RAM[2756] = 32'h00000000,
        RAM[2757] = 32'h00000000,
        RAM[2758] = 32'h00000000,
        RAM[2759] = 32'h00000000,
        RAM[2760] = 32'h00000000,
        RAM[2761] = 32'h00000000,
        RAM[2762] = 32'h00000000,
        RAM[2763] = 32'h00000000,
        RAM[2764] = 32'h00000000,
        RAM[2765] = 32'h00000000,
        RAM[2766] = 32'h00000000,
        RAM[2767] = 32'h00000000,
        RAM[2768] = 32'h00000000,
        RAM[2769] = 32'h00000000,
        RAM[2770] = 32'h00000000,
        RAM[2771] = 32'h00000000,
        RAM[2772] = 32'h00000000,
        RAM[2773] = 32'h00000000,
        RAM[2774] = 32'h00000000,
        RAM[2775] = 32'h00000000,
        RAM[2776] = 32'h00000000,
        RAM[2777] = 32'h00000000,
        RAM[2778] = 32'h00000000,
        RAM[2779] = 32'h00000000,
        RAM[2780] = 32'h00000000,
        RAM[2781] = 32'hffffffff,
        RAM[2782] = 32'h00000000,
        RAM[2783] = 32'h00020000,
        RAM[2784] = 32'h00000000,
        RAM[2785] = 32'h00000000,
        RAM[2786] = 32'h00002b7c,
        RAM[2787] = 32'h00002b7c,
        RAM[2788] = 32'h00002b84,
        RAM[2789] = 32'h00002b84,
        RAM[2790] = 32'h00002b8c,
        RAM[2791] = 32'h00002b8c,
        RAM[2792] = 32'h00002b94,
        RAM[2793] = 32'h00002b94,
        RAM[2794] = 32'h00002b9c,
        RAM[2795] = 32'h00002b9c,
        RAM[2796] = 32'h00002ba4,
        RAM[2797] = 32'h00002ba4,
        RAM[2798] = 32'h00002bac,
        RAM[2799] = 32'h00002bac,
        RAM[2800] = 32'h00002bb4,
        RAM[2801] = 32'h00002bb4,
        RAM[2802] = 32'h00002bbc,
        RAM[2803] = 32'h00002bbc,
        RAM[2804] = 32'h00002bc4,
        RAM[2805] = 32'h00002bc4,
        RAM[2806] = 32'h00002bcc,
        RAM[2807] = 32'h00002bcc,
        RAM[2808] = 32'h00002bd4,
        RAM[2809] = 32'h00002bd4,
        RAM[2810] = 32'h00002bdc,
        RAM[2811] = 32'h00002bdc,
        RAM[2812] = 32'h00002be4,
        RAM[2813] = 32'h00002be4,
        RAM[2814] = 32'h00002bec,
        RAM[2815] = 32'h00002bec,
        RAM[2816] = 32'h00002bf4,
        RAM[2817] = 32'h00002bf4,
        RAM[2818] = 32'h00002bfc,
        RAM[2819] = 32'h00002bfc,
        RAM[2820] = 32'h00002c04,
        RAM[2821] = 32'h00002c04,
        RAM[2822] = 32'h00002c0c,
        RAM[2823] = 32'h00002c0c,
        RAM[2824] = 32'h00002c14,
        RAM[2825] = 32'h00002c14,
        RAM[2826] = 32'h00002c1c,
        RAM[2827] = 32'h00002c1c,
        RAM[2828] = 32'h00002c24,
        RAM[2829] = 32'h00002c24,
        RAM[2830] = 32'h00002c2c,
        RAM[2831] = 32'h00002c2c,
        RAM[2832] = 32'h00002c34,
        RAM[2833] = 32'h00002c34,
        RAM[2834] = 32'h00002c3c,
        RAM[2835] = 32'h00002c3c,
        RAM[2836] = 32'h00002c44,
        RAM[2837] = 32'h00002c44,
        RAM[2838] = 32'h00002c4c,
        RAM[2839] = 32'h00002c4c,
        RAM[2840] = 32'h00002c54,
        RAM[2841] = 32'h00002c54,
        RAM[2842] = 32'h00002c5c,
        RAM[2843] = 32'h00002c5c,
        RAM[2844] = 32'h00002c64,
        RAM[2845] = 32'h00002c64,
        RAM[2846] = 32'h00002c6c,
        RAM[2847] = 32'h00002c6c,
        RAM[2848] = 32'h00002c74,
        RAM[2849] = 32'h00002c74,
        RAM[2850] = 32'h00002c7c,
        RAM[2851] = 32'h00002c7c,
        RAM[2852] = 32'h00002c84,
        RAM[2853] = 32'h00002c84,
        RAM[2854] = 32'h00002c8c,
        RAM[2855] = 32'h00002c8c,
        RAM[2856] = 32'h00002c94,
        RAM[2857] = 32'h00002c94,
        RAM[2858] = 32'h00002c9c,
        RAM[2859] = 32'h00002c9c,
        RAM[2860] = 32'h00002ca4,
        RAM[2861] = 32'h00002ca4,
        RAM[2862] = 32'h00002cac,
        RAM[2863] = 32'h00002cac,
        RAM[2864] = 32'h00002cb4,
        RAM[2865] = 32'h00002cb4,
        RAM[2866] = 32'h00002cbc,
        RAM[2867] = 32'h00002cbc,
        RAM[2868] = 32'h00002cc4,
        RAM[2869] = 32'h00002cc4,
        RAM[2870] = 32'h00002ccc,
        RAM[2871] = 32'h00002ccc,
        RAM[2872] = 32'h00002cd4,
        RAM[2873] = 32'h00002cd4,
        RAM[2874] = 32'h00002cdc,
        RAM[2875] = 32'h00002cdc,
        RAM[2876] = 32'h00002ce4,
        RAM[2877] = 32'h00002ce4,
        RAM[2878] = 32'h00002cec,
        RAM[2879] = 32'h00002cec,
        RAM[2880] = 32'h00002cf4,
        RAM[2881] = 32'h00002cf4,
        RAM[2882] = 32'h00002cfc,
        RAM[2883] = 32'h00002cfc,
        RAM[2884] = 32'h00002d04,
        RAM[2885] = 32'h00002d04,
        RAM[2886] = 32'h00002d0c,
        RAM[2887] = 32'h00002d0c,
        RAM[2888] = 32'h00002d14,
        RAM[2889] = 32'h00002d14,
        RAM[2890] = 32'h00002d1c,
        RAM[2891] = 32'h00002d1c,
        RAM[2892] = 32'h00002d24,
        RAM[2893] = 32'h00002d24,
        RAM[2894] = 32'h00002d2c,
        RAM[2895] = 32'h00002d2c,
        RAM[2896] = 32'h00002d34,
        RAM[2897] = 32'h00002d34,
        RAM[2898] = 32'h00002d3c,
        RAM[2899] = 32'h00002d3c,
        RAM[2900] = 32'h00002d44,
        RAM[2901] = 32'h00002d44,
        RAM[2902] = 32'h00002d4c,
        RAM[2903] = 32'h00002d4c,
        RAM[2904] = 32'h00002d54,
        RAM[2905] = 32'h00002d54,
        RAM[2906] = 32'h00002d5c,
        RAM[2907] = 32'h00002d5c,
        RAM[2908] = 32'h00002d64,
        RAM[2909] = 32'h00002d64,
        RAM[2910] = 32'h00002d6c,
        RAM[2911] = 32'h00002d6c,
        RAM[2912] = 32'h00002d74,
        RAM[2913] = 32'h00002d74,
        RAM[2914] = 32'h00002d7c,
        RAM[2915] = 32'h00002d7c,
        RAM[2916] = 32'h00002d84,
        RAM[2917] = 32'h00002d84,
        RAM[2918] = 32'h00002d8c,
        RAM[2919] = 32'h00002d8c,
        RAM[2920] = 32'h00002d94,
        RAM[2921] = 32'h00002d94,
        RAM[2922] = 32'h00002d9c,
        RAM[2923] = 32'h00002d9c,
        RAM[2924] = 32'h00002da4,
        RAM[2925] = 32'h00002da4,
        RAM[2926] = 32'h00002dac,
        RAM[2927] = 32'h00002dac,
        RAM[2928] = 32'h00002db4,
        RAM[2929] = 32'h00002db4,
        RAM[2930] = 32'h00002dbc,
        RAM[2931] = 32'h00002dbc,
        RAM[2932] = 32'h00002dc4,
        RAM[2933] = 32'h00002dc4,
        RAM[2934] = 32'h00002dcc,
        RAM[2935] = 32'h00002dcc,
        RAM[2936] = 32'h00002dd4,
        RAM[2937] = 32'h00002dd4,
        RAM[2938] = 32'h00002ddc,
        RAM[2939] = 32'h00002ddc,
        RAM[2940] = 32'h00002de4,
        RAM[2941] = 32'h00002de4,
        RAM[2942] = 32'h00002dec,
        RAM[2943] = 32'h00002dec,
        RAM[2944] = 32'h00002df4,
        RAM[2945] = 32'h00002df4,
        RAM[2946] = 32'h00002dfc,
        RAM[2947] = 32'h00002dfc,
        RAM[2948] = 32'h00002e04,
        RAM[2949] = 32'h00002e04,
        RAM[2950] = 32'h00002e0c,
        RAM[2951] = 32'h00002e0c,
        RAM[2952] = 32'h00002e14,
        RAM[2953] = 32'h00002e14,
        RAM[2954] = 32'h00002e1c,
        RAM[2955] = 32'h00002e1c,
        RAM[2956] = 32'h00002e24,
        RAM[2957] = 32'h00002e24,
        RAM[2958] = 32'h00002e2c,
        RAM[2959] = 32'h00002e2c,
        RAM[2960] = 32'h00002e34,
        RAM[2961] = 32'h00002e34,
        RAM[2962] = 32'h00002e3c,
        RAM[2963] = 32'h00002e3c,
        RAM[2964] = 32'h00002e44,
        RAM[2965] = 32'h00002e44,
        RAM[2966] = 32'h00002e4c,
        RAM[2967] = 32'h00002e4c,
        RAM[2968] = 32'h00002e54,
        RAM[2969] = 32'h00002e54,
        RAM[2970] = 32'h00002e5c,
        RAM[2971] = 32'h00002e5c,
        RAM[2972] = 32'h00002e64,
        RAM[2973] = 32'h00002e64,
        RAM[2974] = 32'h00002e6c,
        RAM[2975] = 32'h00002e6c,
        RAM[2976] = 32'h00002e74,
        RAM[2977] = 32'h00002e74,
        RAM[2978] = 32'h00002e7c,
        RAM[2979] = 32'h00002e7c,
        RAM[2980] = 32'h00002e84,
        RAM[2981] = 32'h00002e84,
        RAM[2982] = 32'h00002e8c,
        RAM[2983] = 32'h00002e8c,
        RAM[2984] = 32'h00002e94,
        RAM[2985] = 32'h00002e94,
        RAM[2986] = 32'h00002e9c,
        RAM[2987] = 32'h00002e9c,
        RAM[2988] = 32'h00002ea4,
        RAM[2989] = 32'h00002ea4,
        RAM[2990] = 32'h00002eac,
        RAM[2991] = 32'h00002eac,
        RAM[2992] = 32'h00002eb4,
        RAM[2993] = 32'h00002eb4,
        RAM[2994] = 32'h00002ebc,
        RAM[2995] = 32'h00002ebc,
        RAM[2996] = 32'h00002ec4,
        RAM[2997] = 32'h00002ec4,
        RAM[2998] = 32'h00002ecc,
        RAM[2999] = 32'h00002ecc,
        RAM[3000] = 32'h00002ed4,
        RAM[3001] = 32'h00002ed4,
        RAM[3002] = 32'h00002edc,
        RAM[3003] = 32'h00002edc,
        RAM[3004] = 32'h00002ee4,
        RAM[3005] = 32'h00002ee4,
        RAM[3006] = 32'h00002eec,
        RAM[3007] = 32'h00002eec,
        RAM[3008] = 32'h00002ef4,
        RAM[3009] = 32'h00002ef4,
        RAM[3010] = 32'h00002efc,
        RAM[3011] = 32'h00002efc,
        RAM[3012] = 32'h00002f04,
        RAM[3013] = 32'h00002f04,
        RAM[3014] = 32'h00002f0c,
        RAM[3015] = 32'h00002f0c,
        RAM[3016] = 32'h00002f14,
        RAM[3017] = 32'h00002f14,
        RAM[3018] = 32'h00002f1c,
        RAM[3019] = 32'h00002f1c,
        RAM[3020] = 32'h00002f24,
        RAM[3021] = 32'h00002f24,
        RAM[3022] = 32'h00002f2c,
        RAM[3023] = 32'h00002f2c,
        RAM[3024] = 32'h00002f34,
        RAM[3025] = 32'h00002f34,
        RAM[3026] = 32'h00002f3c,
        RAM[3027] = 32'h00002f3c,
        RAM[3028] = 32'h00002f44,
        RAM[3029] = 32'h00002f44,
        RAM[3030] = 32'h00002f4c,
        RAM[3031] = 32'h00002f4c,
        RAM[3032] = 32'h00002f54,
        RAM[3033] = 32'h00002f54,
        RAM[3034] = 32'h00002f5c,
        RAM[3035] = 32'h00002f5c,
        RAM[3036] = 32'h00002f64,
        RAM[3037] = 32'h00002f64,
        RAM[3038] = 32'h00002f6c,
        RAM[3039] = 32'h00002f6c,
        RAM[3040] = 32'h00002f74,
        RAM[3041] = 32'h00002f74,
        RAM[3042] = 32'h00002724,
        RAM[3043] = 32'hffffffff,
        RAM[3044] = 32'h00000000,
        RAM[3045] = 32'hffffffff,
        RAM[3046] = 32'h00000000,
        RAM[3047] = 32'h00000000,
        RAM[3048] = 32'h00000000,
        RAM[3049] = 32'h00000000,
        RAM[3050] = 32'h00000000,
        RAM[3051] = 32'h00000000,
        RAM[3052] = 32'h00000000,
        RAM[3053] = 32'h00000000,
        RAM[3054] = 32'h00000000,
        RAM[3055] = 32'h00000000,
        RAM[3056] = 32'h00000000,
        RAM[3057] = 32'h00000000,
        RAM[3058] = 32'h00000000,
        RAM[3059] = 32'h00000000,
        RAM[3060] = 32'h00000000,
        RAM[3061] = 32'h00000000,
        RAM[3062] = 32'h00000000,
        RAM[3063] = 32'h00000000,
        RAM[3064] = 32'h00000000,
        RAM[3065] = 32'h00000000,
        RAM[3066] = 32'h00000000,
        RAM[3067] = 32'h00000000,
        RAM[3068] = 32'h00000000,
        RAM[3069] = 32'h00000000,
        RAM[3070] = 32'h00000000,
        RAM[3071] = 32'h00000000,
        RAM[3072] = 32'h00000000,
        RAM[3073] = 32'h00000000,
        RAM[3074] = 32'h00000000,
        RAM[3075] = 32'h00000000,
        RAM[3076] = 32'h00000000,
        RAM[3077] = 32'h00000000,
        RAM[3078] = 32'h00000000,
        RAM[3079] = 32'h00000000,
        RAM[3080] = 32'h00000000,
        RAM[3081] = 32'h00000000,
        RAM[3082] = 32'h00000000,
        RAM[3083] = 32'h00000000,
        RAM[3084] = 32'h00000000,
        RAM[3085] = 32'h00000000,
        RAM[3086] = 32'h00000000,
        RAM[3087] = 32'h00000000,
        RAM[3088] = 32'h00000000,
        RAM[3089] = 32'h00000000,
        RAM[3090] = 32'h00000000,
        RAM[3091] = 32'h00000000,
        RAM[3092] = 32'h00000000,
        RAM[3093] = 32'h00000000,
        RAM[3094] = 32'h00000000,
        RAM[3095] = 32'h00000000,
        RAM[3096] = 32'h00000000,
        RAM[3097] = 32'h00000000,
        RAM[3098] = 32'h00000000,
        RAM[3099] = 32'h00000000,
        RAM[3100] = 32'h00000000,
        RAM[3101] = 32'h00000000,
        RAM[3102] = 32'h00000000,
        RAM[3103] = 32'h00000000,
        RAM[3104] = 32'h00000000,
        RAM[3105] = 32'h00000000,
        RAM[3106] = 32'h00000000,
        RAM[3107] = 32'h00000000,
        RAM[3108] = 32'h00000000,
        RAM[3109] = 32'h00000000,
        RAM[3110] = 32'h00000000,
        RAM[3111] = 32'h00000000,
        RAM[3112] = 32'h00000000,
        RAM[3113] = 32'h00000000,
        RAM[3114] = 32'h00000000,
        RAM[3115] = 32'h00000000,
        RAM[3116] = 32'h00000000,
        RAM[3117] = 32'h00000000,
        RAM[3118] = 32'h00000000,
        RAM[3119] = 32'h00000000,
        RAM[3120] = 32'h00000000,
        RAM[3121] = 32'h00000000,
        RAM[3122] = 32'h00000000,
        RAM[3123] = 32'h00000000,
        RAM[3124] = 32'h00000000,
        RAM[3125] = 32'h00000000,
        RAM[3126] = 32'h00000000,
        RAM[3127] = 32'h00000000,
        RAM[3128] = 32'h00000000,
        RAM[3129] = 32'h00000000,
        RAM[3130] = 32'h00000000,
        RAM[3131] = 32'h00000000,
        RAM[3132] = 32'h00000000,
        RAM[3133] = 32'h00000000,
        RAM[3134] = 32'h00000000,
        RAM[3135] = 32'h00000000,
        RAM[3136] = 32'h00000000,
        RAM[3137] = 32'h00000000,
        RAM[3138] = 32'h00000000,
        RAM[3139] = 32'h00000000,
        RAM[3140] = 32'h00000000,
        RAM[3141] = 32'h00000000,
        RAM[3142] = 32'h00000000,
        RAM[3143] = 32'h00000000,
        RAM[3144] = 32'h00000000,
        RAM[3145] = 32'h00000000,
        RAM[3146] = 32'h00000000,
        RAM[3147] = 32'h00000000,
        RAM[3148] = 32'h00000000,
        RAM[3149] = 32'h00000000,
        RAM[3150] = 32'h00000000,
        RAM[3151] = 32'h00000000,
        RAM[3152] = 32'h00000000,
        RAM[3153] = 32'h00000000,
        RAM[3154] = 32'h00000000,
        RAM[3155] = 32'h00000000,
        RAM[3156] = 32'h00000000,
        RAM[3157] = 32'h00000000,
        RAM[3158] = 32'h00000000,
        RAM[3159] = 32'h00000000,
        RAM[3160] = 32'h00000000,
        RAM[3161] = 32'h00000000,
        RAM[3162] = 32'h00000000,
        RAM[3163] = 32'h00000000,
        RAM[3164] = 32'h00000000,
        RAM[3165] = 32'h00000000,
        RAM[3166] = 32'h00000000,
        RAM[3167] = 32'h00000000,
        RAM[3168] = 32'h00000000,
        RAM[3169] = 32'h00000000,
        RAM[3170] = 32'h00000000,
        RAM[3171] = 32'h00000000,
        RAM[3172] = 32'h00000000,
        RAM[3173] = 32'h00000000,
        RAM[3174] = 32'h00000000,
        RAM[3175] = 32'h00000000,
        RAM[3176] = 32'h00000000,
        RAM[3177] = 32'h00000000,
        RAM[3178] = 32'h00000000,
        RAM[3179] = 32'h00000000,
        RAM[3180] = 32'h00000000,
        RAM[3181] = 32'h00000000,
        RAM[3182] = 32'h00000000,
        RAM[3183] = 32'h00000000,
        RAM[3184] = 32'h00000000,
        RAM[3185] = 32'h00000000,
        RAM[3186] = 32'h00000000,
        RAM[3187] = 32'h00000000,
        RAM[3188] = 32'h00000000,
        RAM[3189] = 32'h00000000,
        RAM[3190] = 32'h00000000,
        RAM[3191] = 32'h00000000,
        RAM[3192] = 32'h00000000,
        RAM[3193] = 32'h00000000,
        RAM[3194] = 32'h00000000,
        RAM[3195] = 32'h00000000,
        RAM[3196] = 32'h00000000,
        RAM[3197] = 32'h00000000,
        RAM[3198] = 32'h00000000,
        RAM[3199] = 32'h00000000,
        RAM[3200] = 32'h00000000,
        RAM[3201] = 32'h00000000,
        RAM[3202] = 32'h00000000,
        RAM[3203] = 32'h00000000,
        RAM[3204] = 32'h00000000,
        RAM[3205] = 32'h00000000,
        RAM[3206] = 32'h00000000,
        RAM[3207] = 32'h00000000,
        RAM[3208] = 32'h00000000,
        RAM[3209] = 32'h00000000,
        RAM[3210] = 32'h00000000,
        RAM[3211] = 32'h00000000,
        RAM[3212] = 32'h00000000,
        RAM[3213] = 32'h00000000,
        RAM[3214] = 32'h00000000,
        RAM[3215] = 32'h00000000,
        RAM[3216] = 32'h00000000,
        RAM[3217] = 32'h00000000,
        RAM[3218] = 32'h00000000,
        RAM[3219] = 32'h00000000,
        RAM[3220] = 32'h00000000,
        RAM[3221] = 32'h00000000,
        RAM[3222] = 32'h00000000,
        RAM[3223] = 32'h00000000,
        RAM[3224] = 32'h00000000,
        RAM[3225] = 32'h00000000,
        RAM[3226] = 32'h00000000,
        RAM[3227] = 32'h00000000,
        RAM[3228] = 32'h00000000,
        RAM[3229] = 32'h00000000,
        RAM[3230] = 32'h00000000,
        RAM[3231] = 32'h00000000,
        RAM[3232] = 32'h00000000,
        RAM[3233] = 32'h00000000,
        RAM[3234] = 32'h00000000,
        RAM[3235] = 32'h00000000,
        RAM[3236] = 32'h00000000,
        RAM[3237] = 32'h00000000,
        RAM[3238] = 32'h00000000,
        RAM[3239] = 32'h00000000,
        RAM[3240] = 32'h00000000,
        RAM[3241] = 32'h00000000,
        RAM[3242] = 32'h00000000,
        RAM[3243] = 32'h00000000,
        RAM[3244] = 32'h00000000,
        RAM[3245] = 32'h00000000,
        RAM[3246] = 32'h00000000,
        RAM[3247] = 32'h00000000,
        RAM[3248] = 32'h00000000,
        RAM[3249] = 32'h00000000,
        RAM[3250] = 32'h00000000,
        RAM[3251] = 32'h00000000,
        RAM[3252] = 32'h00000000,
        RAM[3253] = 32'h00000000,
        RAM[3254] = 32'h00000000,
        RAM[3255] = 32'h00000000,
        RAM[3256] = 32'h00000000,
        RAM[3257] = 32'h00000000,
        RAM[3258] = 32'h00000000,
        RAM[3259] = 32'h00000000,
        RAM[3260] = 32'h00000000,
        RAM[3261] = 32'h00000000,
        RAM[3262] = 32'h00000000,
        RAM[3263] = 32'h00000000,
        RAM[3264] = 32'h00000000,
        RAM[3265] = 32'h00000000,
        RAM[3266] = 32'h00000000,
        RAM[3267] = 32'h00000000,
        RAM[3268] = 32'h00000000,
        RAM[3269] = 32'h00000000,
        RAM[3270] = 32'h00000000,
        RAM[3271] = 32'h00000000,
        RAM[3272] = 32'h00000000,
        RAM[3273] = 32'h00000000,
        RAM[3274] = 32'h00000000,
        RAM[3275] = 32'h00000000,
        RAM[3276] = 32'h00000000,
        RAM[3277] = 32'h00000000,
        RAM[3278] = 32'h00000000,
        RAM[3279] = 32'h00000000,
        RAM[3280] = 32'h00000000,
        RAM[3281] = 32'h00000000,
        RAM[3282] = 32'h00000000,
        RAM[3283] = 32'h00000000,
        RAM[3284] = 32'h00000000,
        RAM[3285] = 32'h00000000,
        RAM[3286] = 32'h00000000,
        RAM[3287] = 32'h00000000,
        RAM[3288] = 32'h00000000,
        RAM[3289] = 32'h00000000,
        RAM[3290] = 32'h00000000,
        RAM[3291] = 32'h00000000,
        RAM[3292] = 32'h00000000,
        RAM[3293] = 32'h00000000,
        RAM[3294] = 32'h00000000,
        RAM[3295] = 32'h00000000,
        RAM[3296] = 32'h00000000,
        RAM[3297] = 32'h00000000,
        RAM[3298] = 32'h00000000,
        RAM[3299] = 32'h00000000,
        RAM[3300] = 32'h00000000,
        RAM[3301] = 32'h00000000,
        RAM[3302] = 32'h00000000,
        RAM[3303] = 32'h00000000,
        RAM[3304] = 32'h00000000,
        RAM[3305] = 32'h00000000,
        RAM[3306] = 32'h00000000,
        RAM[3307] = 32'h00000000,
        RAM[3308] = 32'h00000000,
        RAM[3309] = 32'h00000000,
        RAM[3310] = 32'h00000000,
        RAM[3311] = 32'h00000000,
        RAM[3312] = 32'h00000000,
        RAM[3313] = 32'h00000000,
        RAM[3314] = 32'h00000000,
        RAM[3315] = 32'h00000000,
        RAM[3316] = 32'h00000000,
        RAM[3317] = 32'h00000000,
        RAM[3318] = 32'h00000000,
        RAM[3319] = 32'h00000000,
        RAM[3320] = 32'h00000000,
        RAM[3321] = 32'h00000000,
        RAM[3322] = 32'h00000000,
        RAM[3323] = 32'h00000000,
        RAM[3324] = 32'h00000000,
        RAM[3325] = 32'h00000000,
        RAM[3326] = 32'h00000000,
        RAM[3327] = 32'h00000000,
        RAM[3328] = 32'h00000000,
        RAM[3329] = 32'h00000000,
        RAM[3330] = 32'h00000000,
        RAM[3331] = 32'h00000000,
        RAM[3332] = 32'h00000000,
        RAM[3333] = 32'h00000000,
        RAM[3334] = 32'h00000000,
        RAM[3335] = 32'h00000000,
        RAM[3336] = 32'h00000000,
        RAM[3337] = 32'h00000000,
        RAM[3338] = 32'h00000000,
        RAM[3339] = 32'h00000000,
        RAM[3340] = 32'h00000000,
        RAM[3341] = 32'h00000000,
        RAM[3342] = 32'h00000000,
        RAM[3343] = 32'h00000000,
        RAM[3344] = 32'h00000000,
        RAM[3345] = 32'h00000000,
        RAM[3346] = 32'h00000000,
        RAM[3347] = 32'h00000000,
        RAM[3348] = 32'h00000000,
        RAM[3349] = 32'h00000000,
        RAM[3350] = 32'h00000000,
        RAM[3351] = 32'h00000000,
        RAM[3352] = 32'h00000000,
        RAM[3353] = 32'h00000000,
        RAM[3354] = 32'h00000000,
        RAM[3355] = 32'h00000000,
        RAM[3356] = 32'h00000000,
        RAM[3357] = 32'h00000000,
        RAM[3358] = 32'h00000000,
        RAM[3359] = 32'h00000000,
        RAM[3360] = 32'h00000000,
        RAM[3361] = 32'h00000000,
        RAM[3362] = 32'h00000000,
        RAM[3363] = 32'h00000000,
        RAM[3364] = 32'h00000000,
        RAM[3365] = 32'h00000000,
        RAM[3366] = 32'h00000000,
        RAM[3367] = 32'h00000000,
        RAM[3368] = 32'h00000000,
        RAM[3369] = 32'h00000000,
        RAM[3370] = 32'h00000000,
        RAM[3371] = 32'h00000000,
        RAM[3372] = 32'h00000000,
        RAM[3373] = 32'h00000000,
        RAM[3374] = 32'h00000000,
        RAM[3375] = 32'h00000000,
        RAM[3376] = 32'h00000000,
        RAM[3377] = 32'h00000000,
        RAM[3378] = 32'h00000000,
        RAM[3379] = 32'h00000000,
        RAM[3380] = 32'h00000000,
        RAM[3381] = 32'h00000000,
        RAM[3382] = 32'h00000000,
        RAM[3383] = 32'h00000000,
        RAM[3384] = 32'h00000000,
        RAM[3385] = 32'h00000000,
        RAM[3386] = 32'h00000000,
        RAM[3387] = 32'h00000000,
        RAM[3388] = 32'h00000000,
        RAM[3389] = 32'h00000000,
        RAM[3390] = 32'h00000000,
        RAM[3391] = 32'h00000000,
        RAM[3392] = 32'h00000000,
        RAM[3393] = 32'h00000000,
        RAM[3394] = 32'h00000000,
        RAM[3395] = 32'h00000000,
        RAM[3396] = 32'h00000000,
        RAM[3397] = 32'h00000000,
        RAM[3398] = 32'h00000000,
        RAM[3399] = 32'h00000000,
        RAM[3400] = 32'h00000000,
        RAM[3401] = 32'h00000000,
        RAM[3402] = 32'h00000000,
        RAM[3403] = 32'h00000000,
        RAM[3404] = 32'h00000000,
        RAM[3405] = 32'h00000000,
        RAM[3406] = 32'h00000000,
        RAM[3407] = 32'h00000000,
        RAM[3408] = 32'h00000000,
        RAM[3409] = 32'h00000000,
        RAM[3410] = 32'h00000000,
        RAM[3411] = 32'h00000000,
        RAM[3412] = 32'h00000000,
        RAM[3413] = 32'h00000000,
        RAM[3414] = 32'h00000000,
        RAM[3415] = 32'h00000000,
        RAM[3416] = 32'h00000000,
        RAM[3417] = 32'h00000000,
        RAM[3418] = 32'h00000000,
        RAM[3419] = 32'h00000000,
        RAM[3420] = 32'h00000000,
        RAM[3421] = 32'h00000000,
        RAM[3422] = 32'h00000000,
        RAM[3423] = 32'h00000000,
        RAM[3424] = 32'h00000000,
        RAM[3425] = 32'h00000000,
        RAM[3426] = 32'h00000000,
        RAM[3427] = 32'h00000000,
        RAM[3428] = 32'h00000000,
        RAM[3429] = 32'h00000000,
        RAM[3430] = 32'h00000000,
        RAM[3431] = 32'h00000000,
        RAM[3432] = 32'h00000000,
        RAM[3433] = 32'h00000000,
        RAM[3434] = 32'h00000000,
        RAM[3435] = 32'h00000000,
        RAM[3436] = 32'h00000000,
        RAM[3437] = 32'h00000000,
        RAM[3438] = 32'h00000000,
        RAM[3439] = 32'h00000000,
        RAM[3440] = 32'h00000000,
        RAM[3441] = 32'h00000000,
        RAM[3442] = 32'h00000000,
        RAM[3443] = 32'h00000000,
        RAM[3444] = 32'h00000000,
        RAM[3445] = 32'h00000000,
        RAM[3446] = 32'h00000000,
        RAM[3447] = 32'h00000000,
        RAM[3448] = 32'h00000000,
        RAM[3449] = 32'h00000000,
        RAM[3450] = 32'h00000000,
        RAM[3451] = 32'h00000000,
        RAM[3452] = 32'h00000000,
        RAM[3453] = 32'h00000000,
        RAM[3454] = 32'h00000000,
        RAM[3455] = 32'h00000000,
        RAM[3456] = 32'h00000000,
        RAM[3457] = 32'h00000000,
        RAM[3458] = 32'h00000000,
        RAM[3459] = 32'h00000000,
        RAM[3460] = 32'h00000000,
        RAM[3461] = 32'h00000000,
        RAM[3462] = 32'h00000000,
        RAM[3463] = 32'h00000000,
        RAM[3464] = 32'h00000000,
        RAM[3465] = 32'h00000000,
        RAM[3466] = 32'h00000000,
        RAM[3467] = 32'h00000000,
        RAM[3468] = 32'h00000000,
        RAM[3469] = 32'h00000000,
        RAM[3470] = 32'h00000000,
        RAM[3471] = 32'h00000000,
        RAM[3472] = 32'h00000000,
        RAM[3473] = 32'h00000000,
        RAM[3474] = 32'h00000000,
        RAM[3475] = 32'h00000000,
        RAM[3476] = 32'h00000000,
        RAM[3477] = 32'h00000000,
        RAM[3478] = 32'h00000000,
        RAM[3479] = 32'h00000000,
        RAM[3480] = 32'h00000000,
        RAM[3481] = 32'h00000000,
        RAM[3482] = 32'h00000000,
        RAM[3483] = 32'h00000000,
        RAM[3484] = 32'h00000000,
        RAM[3485] = 32'h00000000,
        RAM[3486] = 32'h00000000,
        RAM[3487] = 32'h00000000,
        RAM[3488] = 32'h00000000,
        RAM[3489] = 32'h00000000,
        RAM[3490] = 32'h00000000,
        RAM[3491] = 32'h00000000,
        RAM[3492] = 32'h00000000,
        RAM[3493] = 32'h00000000,
        RAM[3494] = 32'h00000000,
        RAM[3495] = 32'h00000000,
        RAM[3496] = 32'h00000000,
        RAM[3497] = 32'h00000000,
        RAM[3498] = 32'h00000000,
        RAM[3499] = 32'h00000000,
        RAM[3500] = 32'h00000000,
        RAM[3501] = 32'h00000000,
        RAM[3502] = 32'h00000000,
        RAM[3503] = 32'h00000000,
        RAM[3504] = 32'h00000000,
        RAM[3505] = 32'h00000000,
        RAM[3506] = 32'h00000000,
        RAM[3507] = 32'h00000000,
        RAM[3508] = 32'h00000000,
        RAM[3509] = 32'h00000000,
        RAM[3510] = 32'h00000000,
        RAM[3511] = 32'h00000000,
        RAM[3512] = 32'h00000000,
        RAM[3513] = 32'h00000000,
        RAM[3514] = 32'h00000000,
        RAM[3515] = 32'h00000000,
        RAM[3516] = 32'h00000000,
        RAM[3517] = 32'h00000000,
        RAM[3518] = 32'h00000000,
        RAM[3519] = 32'h00000000,
        RAM[3520] = 32'h00000000,
        RAM[3521] = 32'h00000000,
        RAM[3522] = 32'h00000000,
        RAM[3523] = 32'h00000000,
        RAM[3524] = 32'h00000000,
        RAM[3525] = 32'h00000000,
        RAM[3526] = 32'h00000000,
        RAM[3527] = 32'h00000000,
        RAM[3528] = 32'h00000000,
        RAM[3529] = 32'h00000000,
        RAM[3530] = 32'h00000000,
        RAM[3531] = 32'h00000000,
        RAM[3532] = 32'h00000000,
        RAM[3533] = 32'h00000000,
        RAM[3534] = 32'h00000000,
        RAM[3535] = 32'h00000000,
        RAM[3536] = 32'h00000000,
        RAM[3537] = 32'h00000000,
        RAM[3538] = 32'h00000000,
        RAM[3539] = 32'h00000000,
        RAM[3540] = 32'h00000000,
        RAM[3541] = 32'h00000000,
        RAM[3542] = 32'h00000000,
        RAM[3543] = 32'h00000000,
        RAM[3544] = 32'h00000000,
        RAM[3545] = 32'h00000000,
        RAM[3546] = 32'h00000000,
        RAM[3547] = 32'h00000000,
        RAM[3548] = 32'h00000000,
        RAM[3549] = 32'h00000000,
        RAM[3550] = 32'h00000000,
        RAM[3551] = 32'h00000000,
        RAM[3552] = 32'h00000000,
        RAM[3553] = 32'h00000000,
        RAM[3554] = 32'h00000000,
        RAM[3555] = 32'h00000000,
        RAM[3556] = 32'h00000000,
        RAM[3557] = 32'h00000000,
        RAM[3558] = 32'h00000000,
        RAM[3559] = 32'h00000000,
        RAM[3560] = 32'h00000000,
        RAM[3561] = 32'h00000000,
        RAM[3562] = 32'h00000000,
        RAM[3563] = 32'h00000000,
        RAM[3564] = 32'h00000000,
        RAM[3565] = 32'h00000000,
        RAM[3566] = 32'h00000000,
        RAM[3567] = 32'h00000000,
        RAM[3568] = 32'h00000000,
        RAM[3569] = 32'h00000000,
        RAM[3570] = 32'h00000000,
        RAM[3571] = 32'h00000000,
        RAM[3572] = 32'h00000000,
        RAM[3573] = 32'h00000000,
        RAM[3574] = 32'h00000000,
        RAM[3575] = 32'h00000000,
        RAM[3576] = 32'h00000000,
        RAM[3577] = 32'h00000000,
        RAM[3578] = 32'h00000000,
        RAM[3579] = 32'h00000000,
        RAM[3580] = 32'h00000000,
        RAM[3581] = 32'h00000000,
        RAM[3582] = 32'h00000000,
        RAM[3583] = 32'h00000000,
        RAM[3584] = 32'h00000000,
        RAM[3585] = 32'h00000000,
        RAM[3586] = 32'h00000000,
        RAM[3587] = 32'h00000000,
        RAM[3588] = 32'h00000000,
        RAM[3589] = 32'h00000000,
        RAM[3590] = 32'h00000000,
        RAM[3591] = 32'h00000000,
        RAM[3592] = 32'h00000000,
        RAM[3593] = 32'h00000000,
        RAM[3594] = 32'h00000000,
        RAM[3595] = 32'h00000000,
        RAM[3596] = 32'h00000000,
        RAM[3597] = 32'h00000000,
        RAM[3598] = 32'h00000000,
        RAM[3599] = 32'h00000000,
        RAM[3600] = 32'h00000000,
        RAM[3601] = 32'h00000000,
        RAM[3602] = 32'h00000000,
        RAM[3603] = 32'h00000000,
        RAM[3604] = 32'h00000000,
        RAM[3605] = 32'h00000000,
        RAM[3606] = 32'h00000000,
        RAM[3607] = 32'h00000000,
        RAM[3608] = 32'h00000000,
        RAM[3609] = 32'h00000000,
        RAM[3610] = 32'h00000000,
        RAM[3611] = 32'h00000000,
        RAM[3612] = 32'h00000000,
        RAM[3613] = 32'h00000000,
        RAM[3614] = 32'h00000000,
        RAM[3615] = 32'h00000000,
        RAM[3616] = 32'h00000000,
        RAM[3617] = 32'h00000000,
        RAM[3618] = 32'h00000000,
        RAM[3619] = 32'h00000000,
        RAM[3620] = 32'h00000000,
        RAM[3621] = 32'h00000000,
        RAM[3622] = 32'h00000000,
        RAM[3623] = 32'h00000000,
        RAM[3624] = 32'h00000000,
        RAM[3625] = 32'h00000000,
        RAM[3626] = 32'h00000000,
        RAM[3627] = 32'h00000000,
        RAM[3628] = 32'h00000000,
        RAM[3629] = 32'h00000000,
        RAM[3630] = 32'h00000000,
        RAM[3631] = 32'h00000000,
        RAM[3632] = 32'h00000000,
        RAM[3633] = 32'h00000000,
        RAM[3634] = 32'h00000000,
        RAM[3635] = 32'h00000000,
        RAM[3636] = 32'h00000000,
        RAM[3637] = 32'h00000000,
        RAM[3638] = 32'h00000000,
        RAM[3639] = 32'h00000000,
        RAM[3640] = 32'h00000000,
        RAM[3641] = 32'h00000000,
        RAM[3642] = 32'h00000000,
        RAM[3643] = 32'h00000000,
        RAM[3644] = 32'h00000000,
        RAM[3645] = 32'h00000000,
        RAM[3646] = 32'h00000000,
        RAM[3647] = 32'h00000000,
        RAM[3648] = 32'h00000000,
        RAM[3649] = 32'h00000000,
        RAM[3650] = 32'h00000000,
        RAM[3651] = 32'h00000000,
        RAM[3652] = 32'h00000000,
        RAM[3653] = 32'h00000000,
        RAM[3654] = 32'h00000000,
        RAM[3655] = 32'h00000000,
        RAM[3656] = 32'h00000000,
        RAM[3657] = 32'h00000000,
        RAM[3658] = 32'h00000000,
        RAM[3659] = 32'h00000000,
        RAM[3660] = 32'h00000000,
        RAM[3661] = 32'h00000000,
        RAM[3662] = 32'h00000000,
        RAM[3663] = 32'h00000000,
        RAM[3664] = 32'h00000000,
        RAM[3665] = 32'h00000000,
        RAM[3666] = 32'h00000000,
        RAM[3667] = 32'h00000000,
        RAM[3668] = 32'h00000000,
        RAM[3669] = 32'h00000000,
        RAM[3670] = 32'h00000000,
        RAM[3671] = 32'h00000000,
        RAM[3672] = 32'h00000000,
        RAM[3673] = 32'h00000000,
        RAM[3674] = 32'h00000000,
        RAM[3675] = 32'h00000000,
        RAM[3676] = 32'h00000000,
        RAM[3677] = 32'h00000000,
        RAM[3678] = 32'h00000000,
        RAM[3679] = 32'h00000000,
        RAM[3680] = 32'h00000000,
        RAM[3681] = 32'h00000000,
        RAM[3682] = 32'h00000000,
        RAM[3683] = 32'h00000000,
        RAM[3684] = 32'h00000000,
        RAM[3685] = 32'h00000000,
        RAM[3686] = 32'h00000000,
        RAM[3687] = 32'h00000000,
        RAM[3688] = 32'h00000000,
        RAM[3689] = 32'h00000000,
        RAM[3690] = 32'h00000000,
        RAM[3691] = 32'h00000000,
        RAM[3692] = 32'h00000000,
        RAM[3693] = 32'h00000000,
        RAM[3694] = 32'h00000000,
        RAM[3695] = 32'h00000000,
        RAM[3696] = 32'h00000000,
        RAM[3697] = 32'h00000000,
        RAM[3698] = 32'h00000000,
        RAM[3699] = 32'h00000000,
        RAM[3700] = 32'h00000000,
        RAM[3701] = 32'h00000000,
        RAM[3702] = 32'h00000000,
        RAM[3703] = 32'h00000000,
        RAM[3704] = 32'h00000000,
        RAM[3705] = 32'h00000000,
        RAM[3706] = 32'h00000000,
        RAM[3707] = 32'h00000000,
        RAM[3708] = 32'h00000000,
        RAM[3709] = 32'h00000000,
        RAM[3710] = 32'h00000000,
        RAM[3711] = 32'h00000000,
        RAM[3712] = 32'h00000000,
        RAM[3713] = 32'h00000000,
        RAM[3714] = 32'h00000000,
        RAM[3715] = 32'h00000000,
        RAM[3716] = 32'h00000000,
        RAM[3717] = 32'h00000000,
        RAM[3718] = 32'h00000000,
        RAM[3719] = 32'h00000000,
        RAM[3720] = 32'h00000000,
        RAM[3721] = 32'h00000000,
        RAM[3722] = 32'h00000000,
        RAM[3723] = 32'h00000000,
        RAM[3724] = 32'h00000000,
        RAM[3725] = 32'h00000000,
        RAM[3726] = 32'h00000000,
        RAM[3727] = 32'h00000000,
        RAM[3728] = 32'h00000000,
        RAM[3729] = 32'h00000000,
        RAM[3730] = 32'h00000000,
        RAM[3731] = 32'h00000000,
        RAM[3732] = 32'h00000000,
        RAM[3733] = 32'h00000000,
        RAM[3734] = 32'h00000000,
        RAM[3735] = 32'h00000000,
        RAM[3736] = 32'h00000000,
        RAM[3737] = 32'h00000000,
        RAM[3738] = 32'h00000000,
        RAM[3739] = 32'h00000000,
        RAM[3740] = 32'h00000000,
        RAM[3741] = 32'h00000000,
        RAM[3742] = 32'h00000000,
        RAM[3743] = 32'h00000000,
        RAM[3744] = 32'h00000000,
        RAM[3745] = 32'h00000000,
        RAM[3746] = 32'h00000000,
        RAM[3747] = 32'h00000000,
        RAM[3748] = 32'h00000000,
        RAM[3749] = 32'h00000000,
        RAM[3750] = 32'h00000000,
        RAM[3751] = 32'h00000000,
        RAM[3752] = 32'h00000000,
        RAM[3753] = 32'h00000000,
        RAM[3754] = 32'h00000000,
        RAM[3755] = 32'h00000000,
        RAM[3756] = 32'h00000000,
        RAM[3757] = 32'h00000000,
        RAM[3758] = 32'h00000000,
        RAM[3759] = 32'h00000000,
        RAM[3760] = 32'h00000000,
        RAM[3761] = 32'h00000000,
        RAM[3762] = 32'h00000000,
        RAM[3763] = 32'h00000000,
        RAM[3764] = 32'h00000000,
        RAM[3765] = 32'h00000000,
        RAM[3766] = 32'h00000000,
        RAM[3767] = 32'h00000000,
        RAM[3768] = 32'h00000000,
        RAM[3769] = 32'h00000000,
        RAM[3770] = 32'h00000000,
        RAM[3771] = 32'h00000000,
        RAM[3772] = 32'h00000000,
        RAM[3773] = 32'h00000000,
        RAM[3774] = 32'h00000000,
        RAM[3775] = 32'h00000000,
        RAM[3776] = 32'h00000000,
        RAM[3777] = 32'h00000000,
        RAM[3778] = 32'h00000000,
        RAM[3779] = 32'h00000000,
        RAM[3780] = 32'h00000000,
        RAM[3781] = 32'h00000000,
        RAM[3782] = 32'h00000000,
        RAM[3783] = 32'h00000000,
        RAM[3784] = 32'h00000000,
        RAM[3785] = 32'h00000000,
        RAM[3786] = 32'h00000000,
        RAM[3787] = 32'h00000000,
        RAM[3788] = 32'h00000000,
        RAM[3789] = 32'h00000000,
        RAM[3790] = 32'h00000000,
        RAM[3791] = 32'h00000000,
        RAM[3792] = 32'h00000000,
        RAM[3793] = 32'h00000000,
        RAM[3794] = 32'h00000000,
        RAM[3795] = 32'h00000000,
        RAM[3796] = 32'h00000000,
        RAM[3797] = 32'h00000000,
        RAM[3798] = 32'h00000000,
        RAM[3799] = 32'h00000000,
        RAM[3800] = 32'h00000000,
        RAM[3801] = 32'h00000000,
        RAM[3802] = 32'h00000000,
        RAM[3803] = 32'h00000000,
        RAM[3804] = 32'h00000000,
        RAM[3805] = 32'h00000000,
        RAM[3806] = 32'h00000000,
        RAM[3807] = 32'h00000000,
        RAM[3808] = 32'h00000000,
        RAM[3809] = 32'h00000000,
        RAM[3810] = 32'h00000000,
        RAM[3811] = 32'h00000000,
        RAM[3812] = 32'h00000000,
        RAM[3813] = 32'h00000000,
        RAM[3814] = 32'h00000000,
        RAM[3815] = 32'h00000000,
        RAM[3816] = 32'h00000000,
        RAM[3817] = 32'h00000000,
        RAM[3818] = 32'h00000000,
        RAM[3819] = 32'h00000000,
        RAM[3820] = 32'h00000000,
        RAM[3821] = 32'h00000000,
        RAM[3822] = 32'h00000000,
        RAM[3823] = 32'h00000000,
        RAM[3824] = 32'h00000000,
        RAM[3825] = 32'h00000000,
        RAM[3826] = 32'h00000000,
        RAM[3827] = 32'h00000000,
        RAM[3828] = 32'h00000000,
        RAM[3829] = 32'h00000000,
        RAM[3830] = 32'h00000000,
        RAM[3831] = 32'h00000000,
        RAM[3832] = 32'h00000000,
        RAM[3833] = 32'h00000000,
        RAM[3834] = 32'h00000000,
        RAM[3835] = 32'h00000000,
        RAM[3836] = 32'h00000000,
        RAM[3837] = 32'h00000000,
        RAM[3838] = 32'h00000000,
        RAM[3839] = 32'h00000000,
        RAM[3840] = 32'h00000000,
        RAM[3841] = 32'h00000000,
        RAM[3842] = 32'h00000000,
        RAM[3843] = 32'h00000000,
        RAM[3844] = 32'h00000000,
        RAM[3845] = 32'h00000000,
        RAM[3846] = 32'h00000000,
        RAM[3847] = 32'h00000000,
        RAM[3848] = 32'h00000000,
        RAM[3849] = 32'h00000000,
        RAM[3850] = 32'h00000000,
        RAM[3851] = 32'h00000000,
        RAM[3852] = 32'h00000000,
        RAM[3853] = 32'h00000000,
        RAM[3854] = 32'h00000000,
        RAM[3855] = 32'h00000000,
        RAM[3856] = 32'h00000000,
        RAM[3857] = 32'h00000000,
        RAM[3858] = 32'h00000000,
        RAM[3859] = 32'h00000000,
        RAM[3860] = 32'h00000000,
        RAM[3861] = 32'h00000000,
        RAM[3862] = 32'h00000000,
        RAM[3863] = 32'h00000000,
        RAM[3864] = 32'h00000000,
        RAM[3865] = 32'h00000000,
        RAM[3866] = 32'h00000000,
        RAM[3867] = 32'h00000000,
        RAM[3868] = 32'h00000000,
        RAM[3869] = 32'h00000000,
        RAM[3870] = 32'h00000000,
        RAM[3871] = 32'h00000000,
        RAM[3872] = 32'h00000000,
        RAM[3873] = 32'h00000000,
        RAM[3874] = 32'h00000000,
        RAM[3875] = 32'h00000000,
        RAM[3876] = 32'h00000000,
        RAM[3877] = 32'h00000000,
        RAM[3878] = 32'h00000000,
        RAM[3879] = 32'h00000000,
        RAM[3880] = 32'h00000000,
        RAM[3881] = 32'h00000000,
        RAM[3882] = 32'h00000000,
        RAM[3883] = 32'h00000000,
        RAM[3884] = 32'h00000000,
        RAM[3885] = 32'h00000000,
        RAM[3886] = 32'h00000000,
        RAM[3887] = 32'h00000000,
        RAM[3888] = 32'h00000000,
        RAM[3889] = 32'h00000000,
        RAM[3890] = 32'h00000000,
        RAM[3891] = 32'h00000000,
        RAM[3892] = 32'h00000000,
        RAM[3893] = 32'h00000000,
        RAM[3894] = 32'h00000000,
        RAM[3895] = 32'h00000000,
        RAM[3896] = 32'h00000000,
        RAM[3897] = 32'h00000000,
        RAM[3898] = 32'h00000000,
        RAM[3899] = 32'h00000000,
        RAM[3900] = 32'h00000000,
        RAM[3901] = 32'h00000000,
        RAM[3902] = 32'h00000000,
        RAM[3903] = 32'h00000000,
        RAM[3904] = 32'h00000000,
        RAM[3905] = 32'h00000000,
        RAM[3906] = 32'h00000000,
        RAM[3907] = 32'h00000000,
        RAM[3908] = 32'h00000000,
        RAM[3909] = 32'h00000000,
        RAM[3910] = 32'h00000000,
        RAM[3911] = 32'h00000000,
        RAM[3912] = 32'h00000000,
        RAM[3913] = 32'h00000000,
        RAM[3914] = 32'h00000000,
        RAM[3915] = 32'h00000000,
        RAM[3916] = 32'h00000000,
        RAM[3917] = 32'h00000000,
        RAM[3918] = 32'h00000000,
        RAM[3919] = 32'h00000000,
        RAM[3920] = 32'h00000000,
        RAM[3921] = 32'h00000000,
        RAM[3922] = 32'h00000000,
        RAM[3923] = 32'h00000000,
        RAM[3924] = 32'h00000000,
        RAM[3925] = 32'h00000000,
        RAM[3926] = 32'h00000000,
        RAM[3927] = 32'h00000000,
        RAM[3928] = 32'h00000000,
        RAM[3929] = 32'h00000000,
        RAM[3930] = 32'h00000000,
        RAM[3931] = 32'h00000000,
        RAM[3932] = 32'h00000000,
        RAM[3933] = 32'h00000000,
        RAM[3934] = 32'h00000000,
        RAM[3935] = 32'h00000000,
        RAM[3936] = 32'h00000000,
        RAM[3937] = 32'h00000000,
        RAM[3938] = 32'h00000000,
        RAM[3939] = 32'h00000000,
        RAM[3940] = 32'h00000000,
        RAM[3941] = 32'h00000000,
        RAM[3942] = 32'h00000000,
        RAM[3943] = 32'h00000000,
        RAM[3944] = 32'h00000000,
        RAM[3945] = 32'h00000000,
        RAM[3946] = 32'h00000000,
        RAM[3947] = 32'h00000000,
        RAM[3948] = 32'h00000000,
        RAM[3949] = 32'h00000000,
        RAM[3950] = 32'h00000000,
        RAM[3951] = 32'h00000000,
        RAM[3952] = 32'h00000000,
        RAM[3953] = 32'h00000000,
        RAM[3954] = 32'h00000000,
        RAM[3955] = 32'h00000000,
        RAM[3956] = 32'h00000000,
        RAM[3957] = 32'h00000000,
        RAM[3958] = 32'h00000000,
        RAM[3959] = 32'h00000000,
        RAM[3960] = 32'h00000000,
        RAM[3961] = 32'h00000000,
        RAM[3962] = 32'h00000000,
        RAM[3963] = 32'h00000000,
        RAM[3964] = 32'h00000000,
        RAM[3965] = 32'h00000000,
        RAM[3966] = 32'h00000000,
        RAM[3967] = 32'h00000000,
        RAM[3968] = 32'h00000000,
        RAM[3969] = 32'h00000000,
        RAM[3970] = 32'h00000000,
        RAM[3971] = 32'h00000000,
        RAM[3972] = 32'h00000000,
        RAM[3973] = 32'h00000000,
        RAM[3974] = 32'h00000000,
        RAM[3975] = 32'h00000000,
        RAM[3976] = 32'h00000000,
        RAM[3977] = 32'h00000000,
        RAM[3978] = 32'h00000000,
        RAM[3979] = 32'h00000000,
        RAM[3980] = 32'h00000000,
        RAM[3981] = 32'h00000000,
        RAM[3982] = 32'h00000000,
        RAM[3983] = 32'h00000000,
        RAM[3984] = 32'h00000000,
        RAM[3985] = 32'h00000000,
        RAM[3986] = 32'h00000000,
        RAM[3987] = 32'h00000000,
        RAM[3988] = 32'h00000000,
        RAM[3989] = 32'h00000000,
        RAM[3990] = 32'h00000000,
        RAM[3991] = 32'h00000000,
        RAM[3992] = 32'h00000000,
        RAM[3993] = 32'h00000000,
        RAM[3994] = 32'h00000000,
        RAM[3995] = 32'h00000000,
        RAM[3996] = 32'h00000000,
        RAM[3997] = 32'h00000000,
        RAM[3998] = 32'h00000000,
        RAM[3999] = 32'h00000000,
        RAM[4000] = 32'h00000000,
        RAM[4001] = 32'h00000000,
        RAM[4002] = 32'h00000000,
        RAM[4003] = 32'h00000000,
        RAM[4004] = 32'h00000000,
        RAM[4005] = 32'h00000000,
        RAM[4006] = 32'h00000000,
        RAM[4007] = 32'h00000000,
        RAM[4008] = 32'h00000000,
        RAM[4009] = 32'h00000000,
        RAM[4010] = 32'h00000000,
        RAM[4011] = 32'h00000000,
        RAM[4012] = 32'h00000000,
        RAM[4013] = 32'h00000000,
        RAM[4014] = 32'h00000000,
        RAM[4015] = 32'h00000000,
        RAM[4016] = 32'h00000000,
        RAM[4017] = 32'h00000000,
        RAM[4018] = 32'h00000000,
        RAM[4019] = 32'h00000000,
        RAM[4020] = 32'h00000000,
        RAM[4021] = 32'h00000000,
        RAM[4022] = 32'h00000000,
        RAM[4023] = 32'h00000000,
        RAM[4024] = 32'h00000000,
        RAM[4025] = 32'h00000000,
        RAM[4026] = 32'h00000000,
        RAM[4027] = 32'h00000000,
        RAM[4028] = 32'h00000000,
        RAM[4029] = 32'h00000000,
        RAM[4030] = 32'h00000000,
        RAM[4031] = 32'h00000000,
        RAM[4032] = 32'h00000000,
        RAM[4033] = 32'h00000000,
        RAM[4034] = 32'h00000000,
        RAM[4035] = 32'h00000000,
        RAM[4036] = 32'h00000000,
        RAM[4037] = 32'h00000000,
        RAM[4038] = 32'h00000000,
        RAM[4039] = 32'h00000000,
        RAM[4040] = 32'h00000000,
        RAM[4041] = 32'h00000000,
        RAM[4042] = 32'h00000000,
        RAM[4043] = 32'h00000000,
        RAM[4044] = 32'h00000000,
        RAM[4045] = 32'h00000000,
        RAM[4046] = 32'h00000000,
        RAM[4047] = 32'h00000000,
        RAM[4048] = 32'h00000000,
        RAM[4049] = 32'h00000000,
        RAM[4050] = 32'h00000000,
        RAM[4051] = 32'h00000000,
        RAM[4052] = 32'h00000000,
        RAM[4053] = 32'h00000000,
        RAM[4054] = 32'h00000000,
        RAM[4055] = 32'h00000000,
        RAM[4056] = 32'h00000000,
        RAM[4057] = 32'h00000000,
        RAM[4058] = 32'h00000000,
        RAM[4059] = 32'h00000000,
        RAM[4060] = 32'h00000000,
        RAM[4061] = 32'h00000000,
        RAM[4062] = 32'h00000000,
        RAM[4063] = 32'h00000000,
        RAM[4064] = 32'h00000000,
        RAM[4065] = 32'h00000000,
        RAM[4066] = 32'h00000000,
        RAM[4067] = 32'h00000000,
        RAM[4068] = 32'h00000000,
        RAM[4069] = 32'h00000000,
        RAM[4070] = 32'h00000000,
        RAM[4071] = 32'h00000000,
        RAM[4072] = 32'h00000000,
        RAM[4073] = 32'h00000000,
        RAM[4074] = 32'h00000000,
        RAM[4075] = 32'h00000000,
        RAM[4076] = 32'h00000000,
        RAM[4077] = 32'h00000000,
        RAM[4078] = 32'h00000000,
        RAM[4079] = 32'h00000000,
        RAM[4080] = 32'h00000000,
        RAM[4081] = 32'h00000000,
        RAM[4082] = 32'h00000000,
        RAM[4083] = 32'h00000000,
        RAM[4084] = 32'h00000000,
        RAM[4085] = 32'h00000000,
        RAM[4086] = 32'h00000000,
        RAM[4087] = 32'h00000000,
        RAM[4088] = 32'h00000000,
        RAM[4089] = 32'h00000000,
        RAM[4090] = 32'h00000000,
        RAM[4091] = 32'h00000000,
        RAM[4092] = 32'h00000000,
        RAM[4093] = 32'h00000000,
        RAM[4094] = 32'h00000000,
        RAM[4095] = 32'h00000000,
        RAM[4096] = 32'h00000000,
        RAM[4097] = 32'h00000000,
        RAM[4098] = 32'h00000000,
        RAM[4099] = 32'h00000000,
        RAM[4100] = 32'h00000000,
        RAM[4101] = 32'h00000000,
        RAM[4102] = 32'h00000000,
        RAM[4103] = 32'h00000000,
        RAM[4104] = 32'h00000000,
        RAM[4105] = 32'h00000000,
        RAM[4106] = 32'h00000000,
        RAM[4107] = 32'h00000000,
        RAM[4108] = 32'h00000000,
        RAM[4109] = 32'h00000000,
        RAM[4110] = 32'h00000000,
        RAM[4111] = 32'h00000000,
        RAM[4112] = 32'h00000000,
        RAM[4113] = 32'h00000000,
        RAM[4114] = 32'h00000000,
        RAM[4115] = 32'h00000000,
        RAM[4116] = 32'h00000000,
        RAM[4117] = 32'h00000000,
        RAM[4118] = 32'h00000000,
        RAM[4119] = 32'h00000000,
        RAM[4120] = 32'h00000000,
        RAM[4121] = 32'h00000000,
        RAM[4122] = 32'h00000000,
        RAM[4123] = 32'h00000000,
        RAM[4124] = 32'h00000000,
        RAM[4125] = 32'h00000000,
        RAM[4126] = 32'h00000000,
        RAM[4127] = 32'h00000000,
        RAM[4128] = 32'h00000000,
        RAM[4129] = 32'h00000000,
        RAM[4130] = 32'h00000000,
        RAM[4131] = 32'h00000000,
        RAM[4132] = 32'h00000000,
        RAM[4133] = 32'h00000000,
        RAM[4134] = 32'h00000000,
        RAM[4135] = 32'h00000000,
        RAM[4136] = 32'h00000000,
        RAM[4137] = 32'h00000000,
        RAM[4138] = 32'h00000000,
        RAM[4139] = 32'h00000000,
        RAM[4140] = 32'h00000000,
        RAM[4141] = 32'h00000000,
        RAM[4142] = 32'h00000000,
        RAM[4143] = 32'h00000000,
        RAM[4144] = 32'h00000000,
        RAM[4145] = 32'h00000000,
        RAM[4146] = 32'h00000000,
        RAM[4147] = 32'h00000000,
        RAM[4148] = 32'h00000000,
        RAM[4149] = 32'h00000000,
        RAM[4150] = 32'h00000000,
        RAM[4151] = 32'h00000000,
        RAM[4152] = 32'h00000000,
        RAM[4153] = 32'h00000000,
        RAM[4154] = 32'h00000000,
        RAM[4155] = 32'h00000000,
        RAM[4156] = 32'h00000000,
        RAM[4157] = 32'h00000000,
        RAM[4158] = 32'h00000000,
        RAM[4159] = 32'h00000000,
        RAM[4160] = 32'h00000000,
        RAM[4161] = 32'h00000000,
        RAM[4162] = 32'h00000000,
        RAM[4163] = 32'h00000000,
        RAM[4164] = 32'h00000000,
        RAM[4165] = 32'h00000000,
        RAM[4166] = 32'h00000000,
        RAM[4167] = 32'h00000000,
        RAM[4168] = 32'h00000000,
        RAM[4169] = 32'h00000000,
        RAM[4170] = 32'h00000000,
        RAM[4171] = 32'h00000000,
        RAM[4172] = 32'h00000000,
        RAM[4173] = 32'h00000000,
        RAM[4174] = 32'h00000000,
        RAM[4175] = 32'h00000000,
        RAM[4176] = 32'h00000000,
        RAM[4177] = 32'h00000000,
        RAM[4178] = 32'h00000000,
        RAM[4179] = 32'h00000000,
        RAM[4180] = 32'h00000000,
        RAM[4181] = 32'h00000000,
        RAM[4182] = 32'h00000000,
        RAM[4183] = 32'h00000000,
        RAM[4184] = 32'h00000000,
        RAM[4185] = 32'h00000000,
        RAM[4186] = 32'h00000000,
        RAM[4187] = 32'h00000000,
        RAM[4188] = 32'h00000000,
        RAM[4189] = 32'h00000000,
        RAM[4190] = 32'h00000000,
        RAM[4191] = 32'h00000000,
        RAM[4192] = 32'h00000000,
        RAM[4193] = 32'h00000000,
        RAM[4194] = 32'h00000000,
        RAM[4195] = 32'h00000000,
        RAM[4196] = 32'h00000000,
        RAM[4197] = 32'h00000000,
        RAM[4198] = 32'h00000000,
        RAM[4199] = 32'h00000000,
        RAM[4200] = 32'h00000000,
        RAM[4201] = 32'h00000000,
        RAM[4202] = 32'h00000000,
        RAM[4203] = 32'h00000000,
        RAM[4204] = 32'h00000000,
        RAM[4205] = 32'h00000000,
        RAM[4206] = 32'h00000000,
        RAM[4207] = 32'h00000000,
        RAM[4208] = 32'h00000000,
        RAM[4209] = 32'h00000000,
        RAM[4210] = 32'h00000000,
        RAM[4211] = 32'h00000000,
        RAM[4212] = 32'h00000000,
        RAM[4213] = 32'h00000000,
        RAM[4214] = 32'h00000000,
        RAM[4215] = 32'h00000000,
        RAM[4216] = 32'h00000000,
        RAM[4217] = 32'h00000000,
        RAM[4218] = 32'h00000000,
        RAM[4219] = 32'h00000000,
        RAM[4220] = 32'h00000000,
        RAM[4221] = 32'h00000000,
        RAM[4222] = 32'h00000000,
        RAM[4223] = 32'h00000000,
        RAM[4224] = 32'h00000000,
        RAM[4225] = 32'h00000000,
        RAM[4226] = 32'h00000000,
        RAM[4227] = 32'h00000000,
        RAM[4228] = 32'h00000000,
        RAM[4229] = 32'h00000000,
        RAM[4230] = 32'h00000000,
        RAM[4231] = 32'h00000000,
        RAM[4232] = 32'h00000000,
        RAM[4233] = 32'h00000000,
        RAM[4234] = 32'h00000000,
        RAM[4235] = 32'h00000000,
        RAM[4236] = 32'h00000000,
        RAM[4237] = 32'h00000000,
        RAM[4238] = 32'h00000000,
        RAM[4239] = 32'h00000000,
        RAM[4240] = 32'h00000000,
        RAM[4241] = 32'h00000000,
        RAM[4242] = 32'h00000000,
        RAM[4243] = 32'h00000000,
        RAM[4244] = 32'h00000000,
        RAM[4245] = 32'h00000000,
        RAM[4246] = 32'h00000000,
        RAM[4247] = 32'h00000000,
        RAM[4248] = 32'h00000000,
        RAM[4249] = 32'h00000000,
        RAM[4250] = 32'h00000000,
        RAM[4251] = 32'h00000000,
        RAM[4252] = 32'h00000000,
        RAM[4253] = 32'h00000000,
        RAM[4254] = 32'h00000000,
        RAM[4255] = 32'h00000000,
        RAM[4256] = 32'h00000000,
        RAM[4257] = 32'h00000000,
        RAM[4258] = 32'h00000000,
        RAM[4259] = 32'h00000000,
        RAM[4260] = 32'h00000000,
        RAM[4261] = 32'h00000000,
        RAM[4262] = 32'h00000000,
        RAM[4263] = 32'h00000000,
        RAM[4264] = 32'h00000000,
        RAM[4265] = 32'h00000000,
        RAM[4266] = 32'h00000000,
        RAM[4267] = 32'h00000000,
        RAM[4268] = 32'h00000000,
        RAM[4269] = 32'h00000000,
        RAM[4270] = 32'h00000000,
        RAM[4271] = 32'h00000000,
        RAM[4272] = 32'h00000000,
        RAM[4273] = 32'h00000000,
        RAM[4274] = 32'h00000000,
        RAM[4275] = 32'h00000000,
        RAM[4276] = 32'h00000000,
        RAM[4277] = 32'h00000000,
        RAM[4278] = 32'h00000000,
        RAM[4279] = 32'h00000000,
        RAM[4280] = 32'h00000000,
        RAM[4281] = 32'h00000000,
        RAM[4282] = 32'h00000000,
        RAM[4283] = 32'h00000000,
        RAM[4284] = 32'h00000000,
        RAM[4285] = 32'h00000000,
        RAM[4286] = 32'h00000000,
        RAM[4287] = 32'h00000000,
        RAM[4288] = 32'h00000000,
        RAM[4289] = 32'h00000000,
        RAM[4290] = 32'h00000000,
        RAM[4291] = 32'h00000000,
        RAM[4292] = 32'h00000000,
        RAM[4293] = 32'h00000000,
        RAM[4294] = 32'h00000000,
        RAM[4295] = 32'h00000000,
        RAM[4296] = 32'h00000000,
        RAM[4297] = 32'h00000000,
        RAM[4298] = 32'h00000000,
        RAM[4299] = 32'h00000000,
        RAM[4300] = 32'h00000000,
        RAM[4301] = 32'h00000000,
        RAM[4302] = 32'h00000000,
        RAM[4303] = 32'h00000000,
        RAM[4304] = 32'h00000000,
        RAM[4305] = 32'h00000000,
        RAM[4306] = 32'h00000000,
        RAM[4307] = 32'h00000000,
        RAM[4308] = 32'h00000000,
        RAM[4309] = 32'h00000000,
        RAM[4310] = 32'h00000000,
        RAM[4311] = 32'h00000000,
        RAM[4312] = 32'h00000000,
        RAM[4313] = 32'h00000000,
        RAM[4314] = 32'h00000000,
        RAM[4315] = 32'h00000000,
        RAM[4316] = 32'h00000000,
        RAM[4317] = 32'h00000000,
        RAM[4318] = 32'h00000000,
        RAM[4319] = 32'h00000000,
        RAM[4320] = 32'h00000000,
        RAM[4321] = 32'h00000000,
        RAM[4322] = 32'h00000000,
        RAM[4323] = 32'h00000000,
        RAM[4324] = 32'h00000000,
        RAM[4325] = 32'h00000000,
        RAM[4326] = 32'h00000000,
        RAM[4327] = 32'h00000000,
        RAM[4328] = 32'h00000000,
        RAM[4329] = 32'h00000000,
        RAM[4330] = 32'h00000000,
        RAM[4331] = 32'h00000000,
        RAM[4332] = 32'h00000000,
        RAM[4333] = 32'h00000000,
        RAM[4334] = 32'h00000000,
        RAM[4335] = 32'h00000000,
        RAM[4336] = 32'h00000000,
        RAM[4337] = 32'h00000000,
        RAM[4338] = 32'h00000000,
        RAM[4339] = 32'h00000000,
        RAM[4340] = 32'h00000000,
        RAM[4341] = 32'h00000000,
        RAM[4342] = 32'h00000000,
        RAM[4343] = 32'h00000000,
        RAM[4344] = 32'h00000000,
        RAM[4345] = 32'h00000000,
        RAM[4346] = 32'h00000000,
        RAM[4347] = 32'h00000000,
        RAM[4348] = 32'h00000000,
        RAM[4349] = 32'h00000000,
        RAM[4350] = 32'h00000000,
        RAM[4351] = 32'h00000000,
        RAM[4352] = 32'h00000000,
        RAM[4353] = 32'h00000000,
        RAM[4354] = 32'h00000000,
        RAM[4355] = 32'h00000000,
        RAM[4356] = 32'h00000000,
        RAM[4357] = 32'h00000000,
        RAM[4358] = 32'h00000000,
        RAM[4359] = 32'h00000000,
        RAM[4360] = 32'h00000000,
        RAM[4361] = 32'h00000000,
        RAM[4362] = 32'h00000000,
        RAM[4363] = 32'h00000000,
        RAM[4364] = 32'h00000000,
        RAM[4365] = 32'h00000000,
        RAM[4366] = 32'h00000000,
        RAM[4367] = 32'h00000000,
        RAM[4368] = 32'h00000000,
        RAM[4369] = 32'h00000000,
        RAM[4370] = 32'h00000000,
        RAM[4371] = 32'h00000000,
        RAM[4372] = 32'h00000000,
        RAM[4373] = 32'h00000000,
        RAM[4374] = 32'h00000000,
        RAM[4375] = 32'h00000000,
        RAM[4376] = 32'h00000000,
        RAM[4377] = 32'h00000000,
        RAM[4378] = 32'h00000000,
        RAM[4379] = 32'h00000000,
        RAM[4380] = 32'h00000000,
        RAM[4381] = 32'h00000000,
        RAM[4382] = 32'h00000000,
        RAM[4383] = 32'h00000000,
        RAM[4384] = 32'h00000000,
        RAM[4385] = 32'h00000000,
        RAM[4386] = 32'h00000000,
        RAM[4387] = 32'h00000000,
        RAM[4388] = 32'h00000000,
        RAM[4389] = 32'h00000000,
        RAM[4390] = 32'h00000000,
        RAM[4391] = 32'h00000000,
        RAM[4392] = 32'h00000000,
        RAM[4393] = 32'h00000000,
        RAM[4394] = 32'h00000000,
        RAM[4395] = 32'h00000000,
        RAM[4396] = 32'h00000000,
        RAM[4397] = 32'h00000000,
        RAM[4398] = 32'h00000000,
        RAM[4399] = 32'h00000000,
        RAM[4400] = 32'h00000000,
        RAM[4401] = 32'h00000000,
        RAM[4402] = 32'h00000000,
        RAM[4403] = 32'h00000000,
        RAM[4404] = 32'h00000000,
        RAM[4405] = 32'h00000000,
        RAM[4406] = 32'h00000000,
        RAM[4407] = 32'h00000000,
        RAM[4408] = 32'h00000000,
        RAM[4409] = 32'h00000000,
        RAM[4410] = 32'h00000000,
        RAM[4411] = 32'h00000000,
        RAM[4412] = 32'h00000000,
        RAM[4413] = 32'h00000000,
        RAM[4414] = 32'h00000000,
        RAM[4415] = 32'h00000000,
        RAM[4416] = 32'h00000000,
        RAM[4417] = 32'h00000000,
        RAM[4418] = 32'h00000000,
        RAM[4419] = 32'h00000000,
        RAM[4420] = 32'h00000000,
        RAM[4421] = 32'h00000000,
        RAM[4422] = 32'h00000000,
        RAM[4423] = 32'h00000000,
        RAM[4424] = 32'h00000000,
        RAM[4425] = 32'h00000000,
        RAM[4426] = 32'h00000000,
        RAM[4427] = 32'h00000000,
        RAM[4428] = 32'h00000000,
        RAM[4429] = 32'h00000000,
        RAM[4430] = 32'h00000000,
        RAM[4431] = 32'h00000000,
        RAM[4432] = 32'h00000000,
        RAM[4433] = 32'h00000000,
        RAM[4434] = 32'h00000000,
        RAM[4435] = 32'h00000000,
        RAM[4436] = 32'h00000000,
        RAM[4437] = 32'h00000000,
        RAM[4438] = 32'h00000000,
        RAM[4439] = 32'h00000000,
        RAM[4440] = 32'h00000000,
        RAM[4441] = 32'h00000000,
        RAM[4442] = 32'h00000000,
        RAM[4443] = 32'h00000000,
        RAM[4444] = 32'h00000000,
        RAM[4445] = 32'h00000000,
        RAM[4446] = 32'h00000000,
        RAM[4447] = 32'h00000000,
        RAM[4448] = 32'h00000000,
        RAM[4449] = 32'h00000000,
        RAM[4450] = 32'h00000000,
        RAM[4451] = 32'h00000000,
        RAM[4452] = 32'h00000000,
        RAM[4453] = 32'h00000000,
        RAM[4454] = 32'h00000000,
        RAM[4455] = 32'h00000000,
        RAM[4456] = 32'h00000000,
        RAM[4457] = 32'h00000000,
        RAM[4458] = 32'h00000000,
        RAM[4459] = 32'h00000000,
        RAM[4460] = 32'h00000000,
        RAM[4461] = 32'h00000000,
        RAM[4462] = 32'h00000000,
        RAM[4463] = 32'h00000000,
        RAM[4464] = 32'h00000000,
        RAM[4465] = 32'h00000000,
        RAM[4466] = 32'h00000000,
        RAM[4467] = 32'h00000000,
        RAM[4468] = 32'h00000000,
        RAM[4469] = 32'h00000000,
        RAM[4470] = 32'h00000000,
        RAM[4471] = 32'h00000000,
        RAM[4472] = 32'h00000000,
        RAM[4473] = 32'h00000000,
        RAM[4474] = 32'h00000000,
        RAM[4475] = 32'h00000000,
        RAM[4476] = 32'h00000000,
        RAM[4477] = 32'h00000000,
        RAM[4478] = 32'h00000000,
        RAM[4479] = 32'h00000000,
        RAM[4480] = 32'h00000000,
        RAM[4481] = 32'h00000000,
        RAM[4482] = 32'h00000000,
        RAM[4483] = 32'h00000000,
        RAM[4484] = 32'h00000000,
        RAM[4485] = 32'h00000000,
        RAM[4486] = 32'h00000000,
        RAM[4487] = 32'h00000000,
        RAM[4488] = 32'h00000000,
        RAM[4489] = 32'h00000000,
        RAM[4490] = 32'h00000000,
        RAM[4491] = 32'h00000000,
        RAM[4492] = 32'h00000000,
        RAM[4493] = 32'h00000000,
        RAM[4494] = 32'h00000000,
        RAM[4495] = 32'h00000000,
        RAM[4496] = 32'h00000000,
        RAM[4497] = 32'h00000000,
        RAM[4498] = 32'h00000000,
        RAM[4499] = 32'h00000000,
        RAM[4500] = 32'h00000000,
        RAM[4501] = 32'h00000000,
        RAM[4502] = 32'h00000000,
        RAM[4503] = 32'h00000000,
        RAM[4504] = 32'h00000000,
        RAM[4505] = 32'h00000000,
        RAM[4506] = 32'h00000000,
        RAM[4507] = 32'h00000000,
        RAM[4508] = 32'h00000000,
        RAM[4509] = 32'h00000000,
        RAM[4510] = 32'h00000000,
        RAM[4511] = 32'h00000000,
        RAM[4512] = 32'h00000000,
        RAM[4513] = 32'h00000000,
        RAM[4514] = 32'h00000000,
        RAM[4515] = 32'h00000000,
        RAM[4516] = 32'h00000000,
        RAM[4517] = 32'h00000000,
        RAM[4518] = 32'h00000000,
        RAM[4519] = 32'h00000000,
        RAM[4520] = 32'h00000000,
        RAM[4521] = 32'h00000000,
        RAM[4522] = 32'h00000000,
        RAM[4523] = 32'h00000000,
        RAM[4524] = 32'h00000000,
        RAM[4525] = 32'h00000000,
        RAM[4526] = 32'h00000000,
        RAM[4527] = 32'h00000000,
        RAM[4528] = 32'h00000000,
        RAM[4529] = 32'h00000000,
        RAM[4530] = 32'h00000000,
        RAM[4531] = 32'h00000000,
        RAM[4532] = 32'h00000000,
        RAM[4533] = 32'h00000000,
        RAM[4534] = 32'h00000000,
        RAM[4535] = 32'h00000000,
        RAM[4536] = 32'h00000000,
        RAM[4537] = 32'h00000000,
        RAM[4538] = 32'h00000000,
        RAM[4539] = 32'h00000000,
        RAM[4540] = 32'h00000000,
        RAM[4541] = 32'h00000000,
        RAM[4542] = 32'h00000000,
        RAM[4543] = 32'h00000000,
        RAM[4544] = 32'h00000000,
        RAM[4545] = 32'h00000000,
        RAM[4546] = 32'h00000000,
        RAM[4547] = 32'h00000000,
        RAM[4548] = 32'h00000000,
        RAM[4549] = 32'h00000000,
        RAM[4550] = 32'h00000000,
        RAM[4551] = 32'h00000000,
        RAM[4552] = 32'h00000000,
        RAM[4553] = 32'h00000000,
        RAM[4554] = 32'h00000000,
        RAM[4555] = 32'h00000000,
        RAM[4556] = 32'h00000000,
        RAM[4557] = 32'h00000000,
        RAM[4558] = 32'h00000000,
        RAM[4559] = 32'h00000000,
        RAM[4560] = 32'h00000000,
        RAM[4561] = 32'h00000000,
        RAM[4562] = 32'h00000000,
        RAM[4563] = 32'h00000000,
        RAM[4564] = 32'h00000000,
        RAM[4565] = 32'h00000000,
        RAM[4566] = 32'h00000000,
        RAM[4567] = 32'h00000000,
        RAM[4568] = 32'h00000000,
        RAM[4569] = 32'h00000000,
        RAM[4570] = 32'h00000000,
        RAM[4571] = 32'h00000000,
        RAM[4572] = 32'h00000000,
        RAM[4573] = 32'h00000000,
        RAM[4574] = 32'h00000000,
        RAM[4575] = 32'h00000000,
        RAM[4576] = 32'h00000000,
        RAM[4577] = 32'h00000000,
        RAM[4578] = 32'h00000000,
        RAM[4579] = 32'h00000000,
        RAM[4580] = 32'h00000000,
        RAM[4581] = 32'h00000000,
        RAM[4582] = 32'h00000000,
        RAM[4583] = 32'h00000000,
        RAM[4584] = 32'h00000000,
        RAM[4585] = 32'h00000000,
        RAM[4586] = 32'h00000000,
        RAM[4587] = 32'h00000000,
        RAM[4588] = 32'h00000000,
        RAM[4589] = 32'h00000000,
        RAM[4590] = 32'h00000000,
        RAM[4591] = 32'h00000000,
        RAM[4592] = 32'h00000000,
        RAM[4593] = 32'h00000000,
        RAM[4594] = 32'h00000000,
        RAM[4595] = 32'h00000000,
        RAM[4596] = 32'h00000000,
        RAM[4597] = 32'h00000000,
        RAM[4598] = 32'h00000000,
        RAM[4599] = 32'h00000000,
        RAM[4600] = 32'h00000000,
        RAM[4601] = 32'h00000000,
        RAM[4602] = 32'h00000000,
        RAM[4603] = 32'h00000000,
        RAM[4604] = 32'h00000000,
        RAM[4605] = 32'h00000000,
        RAM[4606] = 32'h00000000,
        RAM[4607] = 32'h00000000,
        RAM[4608] = 32'h00000000,
        RAM[4609] = 32'h00000000,
        RAM[4610] = 32'h00000000,
        RAM[4611] = 32'h00000000,
        RAM[4612] = 32'h00000000,
        RAM[4613] = 32'h00000000,
        RAM[4614] = 32'h00000000,
        RAM[4615] = 32'h00000000,
        RAM[4616] = 32'h00000000,
        RAM[4617] = 32'h00000000,
        RAM[4618] = 32'h00000000,
        RAM[4619] = 32'h00000000,
        RAM[4620] = 32'h00000000,
        RAM[4621] = 32'h00000000,
        RAM[4622] = 32'h00000000,
        RAM[4623] = 32'h00000000,
        RAM[4624] = 32'h00000000,
        RAM[4625] = 32'h00000000,
        RAM[4626] = 32'h00000000,
        RAM[4627] = 32'h00000000,
        RAM[4628] = 32'h00000000,
        RAM[4629] = 32'h00000000,
        RAM[4630] = 32'h00000000,
        RAM[4631] = 32'h00000000,
        RAM[4632] = 32'h00000000,
        RAM[4633] = 32'h00000000,
        RAM[4634] = 32'h00000000,
        RAM[4635] = 32'h00000000,
        RAM[4636] = 32'h00000000,
        RAM[4637] = 32'h00000000,
        RAM[4638] = 32'h00000000,
        RAM[4639] = 32'h00000000,
        RAM[4640] = 32'h00000000,
        RAM[4641] = 32'h00000000,
        RAM[4642] = 32'h00000000,
        RAM[4643] = 32'h00000000,
        RAM[4644] = 32'h00000000,
        RAM[4645] = 32'h00000000,
        RAM[4646] = 32'h00000000,
        RAM[4647] = 32'h00000000,
        RAM[4648] = 32'h00000000,
        RAM[4649] = 32'h00000000,
        RAM[4650] = 32'h00000000,
        RAM[4651] = 32'h00000000,
        RAM[4652] = 32'h00000000,
        RAM[4653] = 32'h00000000,
        RAM[4654] = 32'h00000000,
        RAM[4655] = 32'h00000000,
        RAM[4656] = 32'h00000000,
        RAM[4657] = 32'h00000000,
        RAM[4658] = 32'h00000000,
        RAM[4659] = 32'h00000000,
        RAM[4660] = 32'h00000000,
        RAM[4661] = 32'h00000000,
        RAM[4662] = 32'h00000000,
        RAM[4663] = 32'h00000000,
        RAM[4664] = 32'h00000000,
        RAM[4665] = 32'h00000000,
        RAM[4666] = 32'h00000000,
        RAM[4667] = 32'h00000000,
        RAM[4668] = 32'h00000000,
        RAM[4669] = 32'h00000000,
        RAM[4670] = 32'h00000000,
        RAM[4671] = 32'h00000000,
        RAM[4672] = 32'h00000000,
        RAM[4673] = 32'h00000000,
        RAM[4674] = 32'h00000000,
        RAM[4675] = 32'h00000000,
        RAM[4676] = 32'h00000000,
        RAM[4677] = 32'h00000000,
        RAM[4678] = 32'h00000000,
        RAM[4679] = 32'h00000000,
        RAM[4680] = 32'h00000000,
        RAM[4681] = 32'h00000000,
        RAM[4682] = 32'h00000000,
        RAM[4683] = 32'h00000000,
        RAM[4684] = 32'h00000000,
        RAM[4685] = 32'h00000000,
        RAM[4686] = 32'h00000000,
        RAM[4687] = 32'h00000000,
        RAM[4688] = 32'h00000000,
        RAM[4689] = 32'h00000000,
        RAM[4690] = 32'h00000000,
        RAM[4691] = 32'h00000000,
        RAM[4692] = 32'h00000000,
        RAM[4693] = 32'h00000000,
        RAM[4694] = 32'h00000000,
        RAM[4695] = 32'h00000000,
        RAM[4696] = 32'h00000000,
        RAM[4697] = 32'h00000000,
        RAM[4698] = 32'h00000000,
        RAM[4699] = 32'h00000000,
        RAM[4700] = 32'h00000000,
        RAM[4701] = 32'h00000000,
        RAM[4702] = 32'h00000000,
        RAM[4703] = 32'h00000000,
        RAM[4704] = 32'h00000000,
        RAM[4705] = 32'h00000000,
        RAM[4706] = 32'h00000000,
        RAM[4707] = 32'h00000000,
        RAM[4708] = 32'h00000000,
        RAM[4709] = 32'h00000000,
        RAM[4710] = 32'h00000000,
        RAM[4711] = 32'h00000000,
        RAM[4712] = 32'h00000000,
        RAM[4713] = 32'h00000000,
        RAM[4714] = 32'h00000000,
        RAM[4715] = 32'h00000000,
        RAM[4716] = 32'h00000000,
        RAM[4717] = 32'h00000000,
        RAM[4718] = 32'h00000000,
        RAM[4719] = 32'h00000000,
        RAM[4720] = 32'h00000000,
        RAM[4721] = 32'h00000000,
        RAM[4722] = 32'h00000000,
        RAM[4723] = 32'h00000000,
        RAM[4724] = 32'h00000000,
        RAM[4725] = 32'h00000000,
        RAM[4726] = 32'h00000000,
        RAM[4727] = 32'h00000000,
        RAM[4728] = 32'h00000000,
        RAM[4729] = 32'h00000000,
        RAM[4730] = 32'h00000000,
        RAM[4731] = 32'h00000000,
        RAM[4732] = 32'h00000000,
        RAM[4733] = 32'h00000000,
        RAM[4734] = 32'h00000000,
        RAM[4735] = 32'h00000000,
        RAM[4736] = 32'h00000000,
        RAM[4737] = 32'h00000000,
        RAM[4738] = 32'h00000000,
        RAM[4739] = 32'h00000000,
        RAM[4740] = 32'h00000000,
        RAM[4741] = 32'h00000000,
        RAM[4742] = 32'h00000000,
        RAM[4743] = 32'h00000000,
        RAM[4744] = 32'h00000000,
        RAM[4745] = 32'h00000000,
        RAM[4746] = 32'h00000000,
        RAM[4747] = 32'h00000000,
        RAM[4748] = 32'h00000000,
        RAM[4749] = 32'h00000000,
        RAM[4750] = 32'h00000000,
        RAM[4751] = 32'h00000000,
        RAM[4752] = 32'h00000000,
        RAM[4753] = 32'h00000000,
        RAM[4754] = 32'h00000000,
        RAM[4755] = 32'h00000000,
        RAM[4756] = 32'h00000000,
        RAM[4757] = 32'h00000000,
        RAM[4758] = 32'h00000000,
        RAM[4759] = 32'h00000000,
        RAM[4760] = 32'h00000000,
        RAM[4761] = 32'h00000000,
        RAM[4762] = 32'h00000000,
        RAM[4763] = 32'h00000000,
        RAM[4764] = 32'h00000000,
        RAM[4765] = 32'h00000000,
        RAM[4766] = 32'h00000000,
        RAM[4767] = 32'h00000000,
        RAM[4768] = 32'h00000000,
        RAM[4769] = 32'h00000000,
        RAM[4770] = 32'h00000000,
        RAM[4771] = 32'h00000000,
        RAM[4772] = 32'h00000000,
        RAM[4773] = 32'h00000000,
        RAM[4774] = 32'h00000000,
        RAM[4775] = 32'h00000000,
        RAM[4776] = 32'h00000000,
        RAM[4777] = 32'h00000000,
        RAM[4778] = 32'h00000000,
        RAM[4779] = 32'h00000000,
        RAM[4780] = 32'h00000000,
        RAM[4781] = 32'h00000000,
        RAM[4782] = 32'h00000000,
        RAM[4783] = 32'h00000000,
        RAM[4784] = 32'h00000000,
        RAM[4785] = 32'h00000000,
        RAM[4786] = 32'h00000000,
        RAM[4787] = 32'h00000000,
        RAM[4788] = 32'h00000000,
        RAM[4789] = 32'h00000000,
        RAM[4790] = 32'h00000000,
        RAM[4791] = 32'h00000000,
        RAM[4792] = 32'h00000000,
        RAM[4793] = 32'h00000000,
        RAM[4794] = 32'h00000000,
        RAM[4795] = 32'h00000000,
        RAM[4796] = 32'h00000000,
        RAM[4797] = 32'h00000000,
        RAM[4798] = 32'h00000000,
        RAM[4799] = 32'h00000000,
        RAM[4800] = 32'h00000000,
        RAM[4801] = 32'h00000000,
        RAM[4802] = 32'h00000000,
        RAM[4803] = 32'h00000000,
        RAM[4804] = 32'h00000000,
        RAM[4805] = 32'h00000000,
        RAM[4806] = 32'h00000000,
        RAM[4807] = 32'h00000000,
        RAM[4808] = 32'h00000000,
        RAM[4809] = 32'h00000000,
        RAM[4810] = 32'h00000000,
        RAM[4811] = 32'h00000000,
        RAM[4812] = 32'h00000000,
        RAM[4813] = 32'h00000000,
        RAM[4814] = 32'h00000000,
        RAM[4815] = 32'h00000000,
        RAM[4816] = 32'h00000000,
        RAM[4817] = 32'h00000000,
        RAM[4818] = 32'h00000000,
        RAM[4819] = 32'h00000000,
        RAM[4820] = 32'h00000000,
        RAM[4821] = 32'h00000000,
        RAM[4822] = 32'h00000000,
        RAM[4823] = 32'h00000000,
        RAM[4824] = 32'h00000000,
        RAM[4825] = 32'h00000000,
        RAM[4826] = 32'h00000000,
        RAM[4827] = 32'h00000000,
        RAM[4828] = 32'h00000000,
        RAM[4829] = 32'h00000000,
        RAM[4830] = 32'h00000000,
        RAM[4831] = 32'h00000000,
        RAM[4832] = 32'h00000000,
        RAM[4833] = 32'h00000000,
        RAM[4834] = 32'h00000000,
        RAM[4835] = 32'h00000000,
        RAM[4836] = 32'h00000000,
        RAM[4837] = 32'h00000000,
        RAM[4838] = 32'h00000000,
        RAM[4839] = 32'h00000000,
        RAM[4840] = 32'h00000000,
        RAM[4841] = 32'h00000000,
        RAM[4842] = 32'h00000000,
        RAM[4843] = 32'h00000000,
        RAM[4844] = 32'h00000000,
        RAM[4845] = 32'h00000000,
        RAM[4846] = 32'h00000000,
        RAM[4847] = 32'h00000000,
        RAM[4848] = 32'h00000000,
        RAM[4849] = 32'h00000000,
        RAM[4850] = 32'h00000000,
        RAM[4851] = 32'h00000000,
        RAM[4852] = 32'h00000000,
        RAM[4853] = 32'h00000000,
        RAM[4854] = 32'h00000000,
        RAM[4855] = 32'h00000000,
        RAM[4856] = 32'h00000000,
        RAM[4857] = 32'h00000000,
        RAM[4858] = 32'h00000000,
        RAM[4859] = 32'h00000000,
        RAM[4860] = 32'h00000000,
        RAM[4861] = 32'h00000000,
        RAM[4862] = 32'h00000000,
        RAM[4863] = 32'h00000000,
        RAM[4864] = 32'h00000000,
        RAM[4865] = 32'h00000000,
        RAM[4866] = 32'h00000000,
        RAM[4867] = 32'h00000000,
        RAM[4868] = 32'h00000000,
        RAM[4869] = 32'h00000000,
        RAM[4870] = 32'h00000000,
        RAM[4871] = 32'h00000000,
        RAM[4872] = 32'h00000000,
        RAM[4873] = 32'h00000000,
        RAM[4874] = 32'h00000000,
        RAM[4875] = 32'h00000000,
        RAM[4876] = 32'h00000000,
        RAM[4877] = 32'h00000000,
        RAM[4878] = 32'h00000000,
        RAM[4879] = 32'h00000000,
        RAM[4880] = 32'h00000000,
        RAM[4881] = 32'h00000000,
        RAM[4882] = 32'h00000000,
        RAM[4883] = 32'h00000000,
        RAM[4884] = 32'h00000000,
        RAM[4885] = 32'h00000000,
        RAM[4886] = 32'h00000000,
        RAM[4887] = 32'h00000000,
        RAM[4888] = 32'h00000000,
        RAM[4889] = 32'h00000000,
        RAM[4890] = 32'h00000000,
        RAM[4891] = 32'h00000000,
        RAM[4892] = 32'h00000000,
        RAM[4893] = 32'h00000000,
        RAM[4894] = 32'h00000000,
        RAM[4895] = 32'h00000000,
        RAM[4896] = 32'h00000000,
        RAM[4897] = 32'h00000000,
        RAM[4898] = 32'h00000000,
        RAM[4899] = 32'h00000000,
        RAM[4900] = 32'h00000000,
        RAM[4901] = 32'h00000000,
        RAM[4902] = 32'h00000000,
        RAM[4903] = 32'h00000000,
        RAM[4904] = 32'h00000000,
        RAM[4905] = 32'h00000000,
        RAM[4906] = 32'h00000000,
        RAM[4907] = 32'h00000000,
        RAM[4908] = 32'h00000000,
        RAM[4909] = 32'h00000000,
        RAM[4910] = 32'h00000000,
        RAM[4911] = 32'h00000000,
        RAM[4912] = 32'h00000000,
        RAM[4913] = 32'h00000000,
        RAM[4914] = 32'h00000000,
        RAM[4915] = 32'h00000000,
        RAM[4916] = 32'h00000000,
        RAM[4917] = 32'h00000000,
        RAM[4918] = 32'h00000000,
        RAM[4919] = 32'h00000000,
        RAM[4920] = 32'h00000000,
        RAM[4921] = 32'h00000000,
        RAM[4922] = 32'h00000000,
        RAM[4923] = 32'h00000000,
        RAM[4924] = 32'h00000000,
        RAM[4925] = 32'h00000000,
        RAM[4926] = 32'h00000000,
        RAM[4927] = 32'h00000000,
        RAM[4928] = 32'h00000000,
        RAM[4929] = 32'h00000000,
        RAM[4930] = 32'h00000000,
        RAM[4931] = 32'h00000000,
        RAM[4932] = 32'h00000000,
        RAM[4933] = 32'h00000000,
        RAM[4934] = 32'h00000000,
        RAM[4935] = 32'h00000000,
        RAM[4936] = 32'h00000000,
        RAM[4937] = 32'h00000000,
        RAM[4938] = 32'h00000000,
        RAM[4939] = 32'h00000000,
        RAM[4940] = 32'h00000000,
        RAM[4941] = 32'h00000000,
        RAM[4942] = 32'h00000000,
        RAM[4943] = 32'h00000000,
        RAM[4944] = 32'h00000000,
        RAM[4945] = 32'h00000000,
        RAM[4946] = 32'h00000000,
        RAM[4947] = 32'h00000000,
        RAM[4948] = 32'h00000000,
        RAM[4949] = 32'h00000000,
        RAM[4950] = 32'h00000000,
        RAM[4951] = 32'h00000000,
        RAM[4952] = 32'h00000000,
        RAM[4953] = 32'h00000000,
        RAM[4954] = 32'h00000000,
        RAM[4955] = 32'h00000000,
        RAM[4956] = 32'h00000000,
        RAM[4957] = 32'h00000000,
        RAM[4958] = 32'h00000000,
        RAM[4959] = 32'h00000000,
        RAM[4960] = 32'h00000000,
        RAM[4961] = 32'h00000000,
        RAM[4962] = 32'h00000000,
        RAM[4963] = 32'h00000000,
        RAM[4964] = 32'h00000000,
        RAM[4965] = 32'h00000000,
        RAM[4966] = 32'h00000000,
        RAM[4967] = 32'h00000000,
        RAM[4968] = 32'h00000000,
        RAM[4969] = 32'h00000000,
        RAM[4970] = 32'h00000000,
        RAM[4971] = 32'h00000000,
        RAM[4972] = 32'h00000000,
        RAM[4973] = 32'h00000000,
        RAM[4974] = 32'h00000000,
        RAM[4975] = 32'h00000000,
        RAM[4976] = 32'h00000000,
        RAM[4977] = 32'h00000000,
        RAM[4978] = 32'h00000000,
        RAM[4979] = 32'h00000000,
        RAM[4980] = 32'h00000000,
        RAM[4981] = 32'h00000000,
        RAM[4982] = 32'h00000000,
        RAM[4983] = 32'h00000000,
        RAM[4984] = 32'h00000000,
        RAM[4985] = 32'h00000000,
        RAM[4986] = 32'h00000000,
        RAM[4987] = 32'h00000000,
        RAM[4988] = 32'h00000000,
        RAM[4989] = 32'h00000000,
        RAM[4990] = 32'h00000000,
        RAM[4991] = 32'h00000000,
        RAM[4992] = 32'h00000000,
        RAM[4993] = 32'h00000000,
        RAM[4994] = 32'h00000000,
        RAM[4995] = 32'h00000000,
        RAM[4996] = 32'h00000000,
        RAM[4997] = 32'h00000000,
        RAM[4998] = 32'h00000000,
        RAM[4999] = 32'h00000000,
        RAM[5000] = 32'h00000000,
        RAM[5001] = 32'h00000000,
        RAM[5002] = 32'h00000000,
        RAM[5003] = 32'h00000000,
        RAM[5004] = 32'h00000000,
        RAM[5005] = 32'h00000000,
        RAM[5006] = 32'h00000000,
        RAM[5007] = 32'h00000000,
        RAM[5008] = 32'h00000000,
        RAM[5009] = 32'h00000000,
        RAM[5010] = 32'h00000000,
        RAM[5011] = 32'h00000000,
        RAM[5012] = 32'h00000000,
        RAM[5013] = 32'h00000000,
        RAM[5014] = 32'h00000000,
        RAM[5015] = 32'h00000000,
        RAM[5016] = 32'h00000000,
        RAM[5017] = 32'h00000000,
        RAM[5018] = 32'h00000000,
        RAM[5019] = 32'h00000000,
        RAM[5020] = 32'h00000000,
        RAM[5021] = 32'h00000000,
        RAM[5022] = 32'h00000000,
        RAM[5023] = 32'h00000000,
        RAM[5024] = 32'h00000000,
        RAM[5025] = 32'h00000000,
        RAM[5026] = 32'h00000000,
        RAM[5027] = 32'h00000000,
        RAM[5028] = 32'h00000000,
        RAM[5029] = 32'h00000000,
        RAM[5030] = 32'h00000000,
        RAM[5031] = 32'h00000000,
        RAM[5032] = 32'h00000000,
        RAM[5033] = 32'h00000000,
        RAM[5034] = 32'h00000000,
        RAM[5035] = 32'h00000000,
        RAM[5036] = 32'h00000000,
        RAM[5037] = 32'h00000000,
        RAM[5038] = 32'h00000000,
        RAM[5039] = 32'h00000000,
        RAM[5040] = 32'h00000000,
        RAM[5041] = 32'h00000000,
        RAM[5042] = 32'h00000000,
        RAM[5043] = 32'h00000000,
        RAM[5044] = 32'h00000000,
        RAM[5045] = 32'h00000000,
        RAM[5046] = 32'h00000000,
        RAM[5047] = 32'h00000000,
        RAM[5048] = 32'h00000000,
        RAM[5049] = 32'h00000000,
        RAM[5050] = 32'h00000000,
        RAM[5051] = 32'h00000000,
        RAM[5052] = 32'h00000000,
        RAM[5053] = 32'h00000000,
        RAM[5054] = 32'h00000000,
        RAM[5055] = 32'h00000000,
        RAM[5056] = 32'h00000000,
        RAM[5057] = 32'h00000000,
        RAM[5058] = 32'h00000000,
        RAM[5059] = 32'h00000000,
        RAM[5060] = 32'h00000000,
        RAM[5061] = 32'h00000000,
        RAM[5062] = 32'h00000000,
        RAM[5063] = 32'h00000000,
        RAM[5064] = 32'h00000000,
        RAM[5065] = 32'h00000000,
        RAM[5066] = 32'h00000000,
        RAM[5067] = 32'h00000000,
        RAM[5068] = 32'h00000000,
        RAM[5069] = 32'h00000000,
        RAM[5070] = 32'h00000000,
        RAM[5071] = 32'h00000000,
        RAM[5072] = 32'h00000000,
        RAM[5073] = 32'h00000000,
        RAM[5074] = 32'h00000000,
        RAM[5075] = 32'h00000000,
        RAM[5076] = 32'h00000000,
        RAM[5077] = 32'h00000000,
        RAM[5078] = 32'h00000000,
        RAM[5079] = 32'h00000000,
        RAM[5080] = 32'h00000000,
        RAM[5081] = 32'h00000000,
        RAM[5082] = 32'h00000000,
        RAM[5083] = 32'h00000000,
        RAM[5084] = 32'h00000000,
        RAM[5085] = 32'h00000000,
        RAM[5086] = 32'h00000000,
        RAM[5087] = 32'h00000000,
        RAM[5088] = 32'h00000000,
        RAM[5089] = 32'h00000000,
        RAM[5090] = 32'h00000000,
        RAM[5091] = 32'h00000000,
        RAM[5092] = 32'h00000000,
        RAM[5093] = 32'h00000000,
        RAM[5094] = 32'h00000000,
        RAM[5095] = 32'h00000000,
        RAM[5096] = 32'h00000000,
        RAM[5097] = 32'h00000000,
        RAM[5098] = 32'h00000000,
        RAM[5099] = 32'h00000000,
        RAM[5100] = 32'h00000000,
        RAM[5101] = 32'h00000000,
        RAM[5102] = 32'h00000000,
        RAM[5103] = 32'h00000000,
        RAM[5104] = 32'h00000000,
        RAM[5105] = 32'h00000000,
        RAM[5106] = 32'h00000000,
        RAM[5107] = 32'h00000000,
        RAM[5108] = 32'h00000000,
        RAM[5109] = 32'h00000000,
        RAM[5110] = 32'h00000000,
        RAM[5111] = 32'h00000000,
        RAM[5112] = 32'h00000000,
        RAM[5113] = 32'h00000000,
        RAM[5114] = 32'h00000000,
        RAM[5115] = 32'h00000000,
        RAM[5116] = 32'h00000000,
        RAM[5117] = 32'h00000000,
        RAM[5118] = 32'h00000000,
        RAM[5119] = 32'h00000000,
        RAM[5120] = 32'h00000000,
        RAM[5121] = 32'h00000000,
        RAM[5122] = 32'h00000000,
        RAM[5123] = 32'h00000000,
        RAM[5124] = 32'h00000000,
        RAM[5125] = 32'h00000000,
        RAM[5126] = 32'h00000000,
        RAM[5127] = 32'h00000000,
        RAM[5128] = 32'h00000000,
        RAM[5129] = 32'h00000000,
        RAM[5130] = 32'h00000000,
        RAM[5131] = 32'h00000000,
        RAM[5132] = 32'h00000000,
        RAM[5133] = 32'h00000000,
        RAM[5134] = 32'h00000000,
        RAM[5135] = 32'h00000000,
        RAM[5136] = 32'h00000000,
        RAM[5137] = 32'h00000000,
        RAM[5138] = 32'h00000000,
        RAM[5139] = 32'h00000000,
        RAM[5140] = 32'h00000000,
        RAM[5141] = 32'h00000000,
        RAM[5142] = 32'h00000000,
        RAM[5143] = 32'h00000000,
        RAM[5144] = 32'h00000000,
        RAM[5145] = 32'h00000000,
        RAM[5146] = 32'h00000000,
        RAM[5147] = 32'h00000000,
        RAM[5148] = 32'h00000000,
        RAM[5149] = 32'h00000000,
        RAM[5150] = 32'h00000000,
        RAM[5151] = 32'h00000000,
        RAM[5152] = 32'h00000000,
        RAM[5153] = 32'h00000000,
        RAM[5154] = 32'h00000000,
        RAM[5155] = 32'h00000000,
        RAM[5156] = 32'h00000000,
        RAM[5157] = 32'h00000000,
        RAM[5158] = 32'h00000000,
        RAM[5159] = 32'h00000000,
        RAM[5160] = 32'h00000000,
        RAM[5161] = 32'h00000000,
        RAM[5162] = 32'h00000000,
        RAM[5163] = 32'h00000000,
        RAM[5164] = 32'h00000000,
        RAM[5165] = 32'h00000000,
        RAM[5166] = 32'h00000000,
        RAM[5167] = 32'h00000000,
        RAM[5168] = 32'h00000000,
        RAM[5169] = 32'h00000000,
        RAM[5170] = 32'h00000000,
        RAM[5171] = 32'h00000000,
        RAM[5172] = 32'h00000000,
        RAM[5173] = 32'h00000000,
        RAM[5174] = 32'h00000000,
        RAM[5175] = 32'h00000000,
        RAM[5176] = 32'h00000000,
        RAM[5177] = 32'h00000000,
        RAM[5178] = 32'h00000000,
        RAM[5179] = 32'h00000000,
        RAM[5180] = 32'h00000000,
        RAM[5181] = 32'h00000000,
        RAM[5182] = 32'h00000000,
        RAM[5183] = 32'h00000000,
        RAM[5184] = 32'h00000000,
        RAM[5185] = 32'h00000000,
        RAM[5186] = 32'h00000000,
        RAM[5187] = 32'h00000000,
        RAM[5188] = 32'h00000000,
        RAM[5189] = 32'h00000000,
        RAM[5190] = 32'h00000000,
        RAM[5191] = 32'h00000000,
        RAM[5192] = 32'h00000000,
        RAM[5193] = 32'h00000000,
        RAM[5194] = 32'h00000000,
        RAM[5195] = 32'h00000000,
        RAM[5196] = 32'h00000000,
        RAM[5197] = 32'h00000000,
        RAM[5198] = 32'h00000000,
        RAM[5199] = 32'h00000000,
        RAM[5200] = 32'h00000000,
        RAM[5201] = 32'h00000000,
        RAM[5202] = 32'h00000000,
        RAM[5203] = 32'h00000000,
        RAM[5204] = 32'h00000000,
        RAM[5205] = 32'h00000000,
        RAM[5206] = 32'h00000000,
        RAM[5207] = 32'h00000000,
        RAM[5208] = 32'h00000000,
        RAM[5209] = 32'h00000000,
        RAM[5210] = 32'h00000000,
        RAM[5211] = 32'h00000000,
        RAM[5212] = 32'h00000000,
        RAM[5213] = 32'h00000000,
        RAM[5214] = 32'h00000000,
        RAM[5215] = 32'h00000000,
        RAM[5216] = 32'h00000000,
        RAM[5217] = 32'h00000000,
        RAM[5218] = 32'h00000000,
        RAM[5219] = 32'h00000000,
        RAM[5220] = 32'h00000000,
        RAM[5221] = 32'h00000000,
        RAM[5222] = 32'h00000000,
        RAM[5223] = 32'h00000000,
        RAM[5224] = 32'h00000000,
        RAM[5225] = 32'h00000000,
        RAM[5226] = 32'h00000000,
        RAM[5227] = 32'h00000000,
        RAM[5228] = 32'h00000000,
        RAM[5229] = 32'h00000000,
        RAM[5230] = 32'h00000000,
        RAM[5231] = 32'h00000000,
        RAM[5232] = 32'h00000000,
        RAM[5233] = 32'h00000000,
        RAM[5234] = 32'h00000000,
        RAM[5235] = 32'h00000000,
        RAM[5236] = 32'h00000000,
        RAM[5237] = 32'h00000000,
        RAM[5238] = 32'h00000000,
        RAM[5239] = 32'h00000000,
        RAM[5240] = 32'h00000000,
        RAM[5241] = 32'h00000000,
        RAM[5242] = 32'h00000000,
        RAM[5243] = 32'h00000000,
        RAM[5244] = 32'h00000000,
        RAM[5245] = 32'h00000000,
        RAM[5246] = 32'h00000000,
        RAM[5247] = 32'h00000000,
        RAM[5248] = 32'h00000000,
        RAM[5249] = 32'h00000000,
        RAM[5250] = 32'h00000000,
        RAM[5251] = 32'h00000000,
        RAM[5252] = 32'h00000000,
        RAM[5253] = 32'h00000000,
        RAM[5254] = 32'h00000000,
        RAM[5255] = 32'h00000000,
        RAM[5256] = 32'h00000000,
        RAM[5257] = 32'h00000000,
        RAM[5258] = 32'h00000000,
        RAM[5259] = 32'h00000000,
        RAM[5260] = 32'h00000000,
        RAM[5261] = 32'h00000000,
        RAM[5262] = 32'h00000000,
        RAM[5263] = 32'h00000000,
        RAM[5264] = 32'h00000000,
        RAM[5265] = 32'h00000000,
        RAM[5266] = 32'h00000000,
        RAM[5267] = 32'h00000000,
        RAM[5268] = 32'h00000000,
        RAM[5269] = 32'h00000000,
        RAM[5270] = 32'h00000000,
        RAM[5271] = 32'h00000000,
        RAM[5272] = 32'h00000000,
        RAM[5273] = 32'h00000000,
        RAM[5274] = 32'h00000000,
        RAM[5275] = 32'h00000000,
        RAM[5276] = 32'h00000000,
        RAM[5277] = 32'h00000000,
        RAM[5278] = 32'h00000000,
        RAM[5279] = 32'h00000000,
        RAM[5280] = 32'h00000000,
        RAM[5281] = 32'h00000000,
        RAM[5282] = 32'h00000000,
        RAM[5283] = 32'h00000000,
        RAM[5284] = 32'h00000000,
        RAM[5285] = 32'h00000000,
        RAM[5286] = 32'h00000000,
        RAM[5287] = 32'h00000000,
        RAM[5288] = 32'h00000000,
        RAM[5289] = 32'h00000000,
        RAM[5290] = 32'h00000000,
        RAM[5291] = 32'h00000000,
        RAM[5292] = 32'h00000000,
        RAM[5293] = 32'h00000000,
        RAM[5294] = 32'h00000000,
        RAM[5295] = 32'h00000000,
        RAM[5296] = 32'h00000000,
        RAM[5297] = 32'h00000000,
        RAM[5298] = 32'h00000000,
        RAM[5299] = 32'h00000000,
        RAM[5300] = 32'h00000000,
        RAM[5301] = 32'h00000000,
        RAM[5302] = 32'h00000000,
        RAM[5303] = 32'h00000000,
        RAM[5304] = 32'h00000000,
        RAM[5305] = 32'h00000000,
        RAM[5306] = 32'h00000000,
        RAM[5307] = 32'h00000000,
        RAM[5308] = 32'h00000000,
        RAM[5309] = 32'h00000000,
        RAM[5310] = 32'h00000000,
        RAM[5311] = 32'h00000000,
        RAM[5312] = 32'h00000000,
        RAM[5313] = 32'h00000000,
        RAM[5314] = 32'h00000000,
        RAM[5315] = 32'h00000000,
        RAM[5316] = 32'h00000000,
        RAM[5317] = 32'h00000000,
        RAM[5318] = 32'h00000000,
        RAM[5319] = 32'h00000000,
        RAM[5320] = 32'h00000000,
        RAM[5321] = 32'h00000000,
        RAM[5322] = 32'h00000000,
        RAM[5323] = 32'h00000000,
        RAM[5324] = 32'h00000000,
        RAM[5325] = 32'h00000000,
        RAM[5326] = 32'h00000000,
        RAM[5327] = 32'h00000000,
        RAM[5328] = 32'h00000000,
        RAM[5329] = 32'h00000000,
        RAM[5330] = 32'h00000000,
        RAM[5331] = 32'h00000000,
        RAM[5332] = 32'h00000000,
        RAM[5333] = 32'h00000000,
        RAM[5334] = 32'h00000000,
        RAM[5335] = 32'h00000000,
        RAM[5336] = 32'h00000000,
        RAM[5337] = 32'h00000000,
        RAM[5338] = 32'h00000000,
        RAM[5339] = 32'h00000000,
        RAM[5340] = 32'h00000000,
        RAM[5341] = 32'h00000000,
        RAM[5342] = 32'h00000000,
        RAM[5343] = 32'h00000000,
        RAM[5344] = 32'h00000000,
        RAM[5345] = 32'h00000000,
        RAM[5346] = 32'h00000000,
        RAM[5347] = 32'h00000000,
        RAM[5348] = 32'h00000000,
        RAM[5349] = 32'h00000000,
        RAM[5350] = 32'h00000000,
        RAM[5351] = 32'h00000000,
        RAM[5352] = 32'h00000000,
        RAM[5353] = 32'h00000000,
        RAM[5354] = 32'h00000000,
        RAM[5355] = 32'h00000000,
        RAM[5356] = 32'h00000000,
        RAM[5357] = 32'h00000000,
        RAM[5358] = 32'h00000000,
        RAM[5359] = 32'h00000000,
        RAM[5360] = 32'h00000000,
        RAM[5361] = 32'h00000000,
        RAM[5362] = 32'h00000000,
        RAM[5363] = 32'h00000000,
        RAM[5364] = 32'h00000000,
        RAM[5365] = 32'h00000000,
        RAM[5366] = 32'h00000000,
        RAM[5367] = 32'h00000000,
        RAM[5368] = 32'h00000000,
        RAM[5369] = 32'h00000000,
        RAM[5370] = 32'h00000000,
        RAM[5371] = 32'h00000000,
        RAM[5372] = 32'h00000000,
        RAM[5373] = 32'h00000000,
        RAM[5374] = 32'h00000000,
        RAM[5375] = 32'h00000000,
        RAM[5376] = 32'h00000000,
        RAM[5377] = 32'h00000000,
        RAM[5378] = 32'h00000000,
        RAM[5379] = 32'h00000000,
        RAM[5380] = 32'h00000000,
        RAM[5381] = 32'h00000000,
        RAM[5382] = 32'h00000000,
        RAM[5383] = 32'h00000000,
        RAM[5384] = 32'h00000000,
        RAM[5385] = 32'h00000000,
        RAM[5386] = 32'h00000000,
        RAM[5387] = 32'h00000000,
        RAM[5388] = 32'h00000000,
        RAM[5389] = 32'h00000000,
        RAM[5390] = 32'h00000000,
        RAM[5391] = 32'h00000000,
        RAM[5392] = 32'h00000000,
        RAM[5393] = 32'h00000000,
        RAM[5394] = 32'h00000000,
        RAM[5395] = 32'h00000000,
        RAM[5396] = 32'h00000000,
        RAM[5397] = 32'h00000000,
        RAM[5398] = 32'h00000000,
        RAM[5399] = 32'h00000000,
        RAM[5400] = 32'h00000000,
        RAM[5401] = 32'h00000000,
        RAM[5402] = 32'h00000000,
        RAM[5403] = 32'h00000000,
        RAM[5404] = 32'h00000000,
        RAM[5405] = 32'h00000000,
        RAM[5406] = 32'h00000000,
        RAM[5407] = 32'h00000000,
        RAM[5408] = 32'h00000000,
        RAM[5409] = 32'h00000000,
        RAM[5410] = 32'h00000000,
        RAM[5411] = 32'h00000000,
        RAM[5412] = 32'h00000000,
        RAM[5413] = 32'h00000000,
        RAM[5414] = 32'h00000000,
        RAM[5415] = 32'h00000000,
        RAM[5416] = 32'h00000000,
        RAM[5417] = 32'h00000000,
        RAM[5418] = 32'h00000000,
        RAM[5419] = 32'h00000000,
        RAM[5420] = 32'h00000000,
        RAM[5421] = 32'h00000000,
        RAM[5422] = 32'h00000000,
        RAM[5423] = 32'h00000000,
        RAM[5424] = 32'h00000000,
        RAM[5425] = 32'h00000000,
        RAM[5426] = 32'h00000000,
        RAM[5427] = 32'h00000000,
        RAM[5428] = 32'h00000000,
        RAM[5429] = 32'h00000000,
        RAM[5430] = 32'h00000000,
        RAM[5431] = 32'h00000000,
        RAM[5432] = 32'h00000000,
        RAM[5433] = 32'h00000000,
        RAM[5434] = 32'h00000000,
        RAM[5435] = 32'h00000000,
        RAM[5436] = 32'h00000000,
        RAM[5437] = 32'h00000000,
        RAM[5438] = 32'h00000000,
        RAM[5439] = 32'h00000000,
        RAM[5440] = 32'h00000000,
        RAM[5441] = 32'h00000000,
        RAM[5442] = 32'h00000000,
        RAM[5443] = 32'h00000000,
        RAM[5444] = 32'h00000000,
        RAM[5445] = 32'h00000000,
        RAM[5446] = 32'h00000000,
        RAM[5447] = 32'h00000000,
        RAM[5448] = 32'h00000000,
        RAM[5449] = 32'h00000000,
        RAM[5450] = 32'h00000000,
        RAM[5451] = 32'h00000000,
        RAM[5452] = 32'h00000000,
        RAM[5453] = 32'h00000000,
        RAM[5454] = 32'h00000000,
        RAM[5455] = 32'h00000000,
        RAM[5456] = 32'h00000000,
        RAM[5457] = 32'h00000000,
        RAM[5458] = 32'h00000000,
        RAM[5459] = 32'h00000000,
        RAM[5460] = 32'h00000000,
        RAM[5461] = 32'h00000000,
        RAM[5462] = 32'h00000000,
        RAM[5463] = 32'h00000000,
        RAM[5464] = 32'h00000000,
        RAM[5465] = 32'h00000000,
        RAM[5466] = 32'h00000000,
        RAM[5467] = 32'h00000000,
        RAM[5468] = 32'h00000000,
        RAM[5469] = 32'h00000000,
        RAM[5470] = 32'h00000000,
        RAM[5471] = 32'h00000000,
        RAM[5472] = 32'h00000000,
        RAM[5473] = 32'h00000000,
        RAM[5474] = 32'h00000000,
        RAM[5475] = 32'h00000000,
        RAM[5476] = 32'h00000000,
        RAM[5477] = 32'h00000000,
        RAM[5478] = 32'h00000000,
        RAM[5479] = 32'h00000000,
        RAM[5480] = 32'h00000000,
        RAM[5481] = 32'h00000000,
        RAM[5482] = 32'h00000000,
        RAM[5483] = 32'h00000000,
        RAM[5484] = 32'h00000000,
        RAM[5485] = 32'h00000000,
        RAM[5486] = 32'h00000000,
        RAM[5487] = 32'h00000000,
        RAM[5488] = 32'h00000000,
        RAM[5489] = 32'h00000000,
        RAM[5490] = 32'h00000000,
        RAM[5491] = 32'h00000000,
        RAM[5492] = 32'h00000000,
        RAM[5493] = 32'h00000000,
        RAM[5494] = 32'h00000000,
        RAM[5495] = 32'h00000000,
        RAM[5496] = 32'h00000000,
        RAM[5497] = 32'h00000000,
        RAM[5498] = 32'h00000000,
        RAM[5499] = 32'h00000000,
        RAM[5500] = 32'h00000000,
        RAM[5501] = 32'h00000000,
        RAM[5502] = 32'h00000000,
        RAM[5503] = 32'h00000000,
        RAM[5504] = 32'h00000000,
        RAM[5505] = 32'h00000000,
        RAM[5506] = 32'h00000000,
        RAM[5507] = 32'h00000000,
        RAM[5508] = 32'h00000000,
        RAM[5509] = 32'h00000000,
        RAM[5510] = 32'h00000000,
        RAM[5511] = 32'h00000000,
        RAM[5512] = 32'h00000000,
        RAM[5513] = 32'h00000000,
        RAM[5514] = 32'h00000000,
        RAM[5515] = 32'h00000000,
        RAM[5516] = 32'h00000000,
        RAM[5517] = 32'h00000000,
        RAM[5518] = 32'h00000000,
        RAM[5519] = 32'h00000000,
        RAM[5520] = 32'h00000000,
        RAM[5521] = 32'h00000000,
        RAM[5522] = 32'h00000000,
        RAM[5523] = 32'h00000000,
        RAM[5524] = 32'h00000000,
        RAM[5525] = 32'h00000000,
        RAM[5526] = 32'h00000000,
        RAM[5527] = 32'h00000000,
        RAM[5528] = 32'h00000000,
        RAM[5529] = 32'h00000000,
        RAM[5530] = 32'h00000000,
        RAM[5531] = 32'h00000000,
        RAM[5532] = 32'h00000000,
        RAM[5533] = 32'h00000000,
        RAM[5534] = 32'h00000000,
        RAM[5535] = 32'h00000000,
        RAM[5536] = 32'h00000000,
        RAM[5537] = 32'h00000000,
        RAM[5538] = 32'h00000000,
        RAM[5539] = 32'h00000000,
        RAM[5540] = 32'h00000000,
        RAM[5541] = 32'h00000000,
        RAM[5542] = 32'h00000000,
        RAM[5543] = 32'h00000000,
        RAM[5544] = 32'h00000000,
        RAM[5545] = 32'h00000000,
        RAM[5546] = 32'h00000000,
        RAM[5547] = 32'h00000000,
        RAM[5548] = 32'h00000000,
        RAM[5549] = 32'h00000000,
        RAM[5550] = 32'h00000000,
        RAM[5551] = 32'h00000000,
        RAM[5552] = 32'h00000000,
        RAM[5553] = 32'h00000000,
        RAM[5554] = 32'h00000000,
        RAM[5555] = 32'h00000000,
        RAM[5556] = 32'h00000000,
        RAM[5557] = 32'h00000000,
        RAM[5558] = 32'h00000000,
        RAM[5559] = 32'h00000000,
        RAM[5560] = 32'h00000000,
        RAM[5561] = 32'h00000000,
        RAM[5562] = 32'h00000000,
        RAM[5563] = 32'h00000000,
        RAM[5564] = 32'h00000000,
        RAM[5565] = 32'h00000000,
        RAM[5566] = 32'h00000000,
        RAM[5567] = 32'h00000000,
        RAM[5568] = 32'h00000000,
        RAM[5569] = 32'h00000000,
        RAM[5570] = 32'h00000000,
        RAM[5571] = 32'h00000000,
        RAM[5572] = 32'h00000000,
        RAM[5573] = 32'h00000000,
        RAM[5574] = 32'h00000000,
        RAM[5575] = 32'h00000000,
        RAM[5576] = 32'h00000000,
        RAM[5577] = 32'h00000000,
        RAM[5578] = 32'h00000000,
        RAM[5579] = 32'h00000000,
        RAM[5580] = 32'h00000000,
        RAM[5581] = 32'h00000000,
        RAM[5582] = 32'h00000000,
        RAM[5583] = 32'h00000000,
        RAM[5584] = 32'h00000000,
        RAM[5585] = 32'h00000000,
        RAM[5586] = 32'h00000000,
        RAM[5587] = 32'h00000000,
        RAM[5588] = 32'h00000000,
        RAM[5589] = 32'h00000000,
        RAM[5590] = 32'h00000000,
        RAM[5591] = 32'h00000000,
        RAM[5592] = 32'h00000000,
        RAM[5593] = 32'h00000000,
        RAM[5594] = 32'h00000000,
        RAM[5595] = 32'h00000000,
        RAM[5596] = 32'h00000000,
        RAM[5597] = 32'h00000000,
        RAM[5598] = 32'h00000000,
        RAM[5599] = 32'h00000000,
        RAM[5600] = 32'h00000000,
        RAM[5601] = 32'h00000000,
        RAM[5602] = 32'h00000000,
        RAM[5603] = 32'h00000000,
        RAM[5604] = 32'h00000000,
        RAM[5605] = 32'h00000000,
        RAM[5606] = 32'h00000000,
        RAM[5607] = 32'h00000000,
        RAM[5608] = 32'h00000000,
        RAM[5609] = 32'h00000000,
        RAM[5610] = 32'h00000000,
        RAM[5611] = 32'h00000000,
        RAM[5612] = 32'h00000000,
        RAM[5613] = 32'h00000000,
        RAM[5614] = 32'h00000000,
        RAM[5615] = 32'h00000000,
        RAM[5616] = 32'h00000000,
        RAM[5617] = 32'h00000000,
        RAM[5618] = 32'h00000000,
        RAM[5619] = 32'h00000000,
        RAM[5620] = 32'h00000000,
        RAM[5621] = 32'h00000000,
        RAM[5622] = 32'h00000000,
        RAM[5623] = 32'h00000000,
        RAM[5624] = 32'h00000000,
        RAM[5625] = 32'h00000000,
        RAM[5626] = 32'h00000000,
        RAM[5627] = 32'h00000000,
        RAM[5628] = 32'h00000000,
        RAM[5629] = 32'h00000000,
        RAM[5630] = 32'h00000000,
        RAM[5631] = 32'h00000000,
        RAM[5632] = 32'h00000000,
        RAM[5633] = 32'h00000000,
        RAM[5634] = 32'h00000000,
        RAM[5635] = 32'h00000000,
        RAM[5636] = 32'h00000000,
        RAM[5637] = 32'h00000000,
        RAM[5638] = 32'h00000000,
        RAM[5639] = 32'h00000000,
        RAM[5640] = 32'h00000000,
        RAM[5641] = 32'h00000000,
        RAM[5642] = 32'h00000000,
        RAM[5643] = 32'h00000000,
        RAM[5644] = 32'h00000000,
        RAM[5645] = 32'h00000000,
        RAM[5646] = 32'h00000000,
        RAM[5647] = 32'h00000000,
        RAM[5648] = 32'h00000000,
        RAM[5649] = 32'h00000000,
        RAM[5650] = 32'h00000000,
        RAM[5651] = 32'h00000000,
        RAM[5652] = 32'h00000000,
        RAM[5653] = 32'h00000000,
        RAM[5654] = 32'h00000000,
        RAM[5655] = 32'h00000000,
        RAM[5656] = 32'h00000000,
        RAM[5657] = 32'h00000000,
        RAM[5658] = 32'h00000000,
        RAM[5659] = 32'h00000000,
        RAM[5660] = 32'h00000000,
        RAM[5661] = 32'h00000000,
        RAM[5662] = 32'h00000000,
        RAM[5663] = 32'h00000000,
        RAM[5664] = 32'h00000000,
        RAM[5665] = 32'h00000000,
        RAM[5666] = 32'h00000000,
        RAM[5667] = 32'h00000000,
        RAM[5668] = 32'h00000000,
        RAM[5669] = 32'h00000000,
        RAM[5670] = 32'h00000000,
        RAM[5671] = 32'h00000000,
        RAM[5672] = 32'h00000000,
        RAM[5673] = 32'h00000000,
        RAM[5674] = 32'h00000000,
        RAM[5675] = 32'h00000000,
        RAM[5676] = 32'h00000000,
        RAM[5677] = 32'h00000000,
        RAM[5678] = 32'h00000000,
        RAM[5679] = 32'h00000000,
        RAM[5680] = 32'h00000000,
        RAM[5681] = 32'h00000000,
        RAM[5682] = 32'h00000000,
        RAM[5683] = 32'h00000000,
        RAM[5684] = 32'h00000000,
        RAM[5685] = 32'h00000000,
        RAM[5686] = 32'h00000000,
        RAM[5687] = 32'h00000000,
        RAM[5688] = 32'h00000000,
        RAM[5689] = 32'h00000000,
        RAM[5690] = 32'h00000000,
        RAM[5691] = 32'h00000000,
        RAM[5692] = 32'h00000000,
        RAM[5693] = 32'h00000000,
        RAM[5694] = 32'h00000000,
        RAM[5695] = 32'h00000000,
        RAM[5696] = 32'h00000000,
        RAM[5697] = 32'h00000000,
        RAM[5698] = 32'h00000000,
        RAM[5699] = 32'h00000000,
        RAM[5700] = 32'h00000000,
        RAM[5701] = 32'h00000000,
        RAM[5702] = 32'h00000000,
        RAM[5703] = 32'h00000000,
        RAM[5704] = 32'h00000000,
        RAM[5705] = 32'h00000000,
        RAM[5706] = 32'h00000000,
        RAM[5707] = 32'h00000000,
        RAM[5708] = 32'h00000000,
        RAM[5709] = 32'h00000000,
        RAM[5710] = 32'h00000000,
        RAM[5711] = 32'h00000000,
        RAM[5712] = 32'h00000000,
        RAM[5713] = 32'h00000000,
        RAM[5714] = 32'h00000000,
        RAM[5715] = 32'h00000000,
        RAM[5716] = 32'h00000000,
        RAM[5717] = 32'h00000000,
        RAM[5718] = 32'h00000000,
        RAM[5719] = 32'h00000000,
        RAM[5720] = 32'h00000000,
        RAM[5721] = 32'h00000000,
        RAM[5722] = 32'h00000000,
        RAM[5723] = 32'h00000000,
        RAM[5724] = 32'h00000000,
        RAM[5725] = 32'h00000000,
        RAM[5726] = 32'h00000000,
        RAM[5727] = 32'h00000000,
        RAM[5728] = 32'h00000000,
        RAM[5729] = 32'h00000000,
        RAM[5730] = 32'h00000000,
        RAM[5731] = 32'h00000000,
        RAM[5732] = 32'h00000000,
        RAM[5733] = 32'h00000000,
        RAM[5734] = 32'h00000000,
        RAM[5735] = 32'h00000000,
        RAM[5736] = 32'h00000000,
        RAM[5737] = 32'h00000000,
        RAM[5738] = 32'h00000000,
        RAM[5739] = 32'h00000000,
        RAM[5740] = 32'h00000000,
        RAM[5741] = 32'h00000000,
        RAM[5742] = 32'h00000000,
        RAM[5743] = 32'h00000000,
        RAM[5744] = 32'h00000000,
        RAM[5745] = 32'h00000000,
        RAM[5746] = 32'h00000000,
        RAM[5747] = 32'h00000000,
        RAM[5748] = 32'h00000000,
        RAM[5749] = 32'h00000000,
        RAM[5750] = 32'h00000000,
        RAM[5751] = 32'h00000000,
        RAM[5752] = 32'h00000000,
        RAM[5753] = 32'h00000000,
        RAM[5754] = 32'h00000000,
        RAM[5755] = 32'h00000000,
        RAM[5756] = 32'h00000000,
        RAM[5757] = 32'h00000000,
        RAM[5758] = 32'h00000000,
        RAM[5759] = 32'h00000000,
        RAM[5760] = 32'h00000000,
        RAM[5761] = 32'h00000000,
        RAM[5762] = 32'h00000000,
        RAM[5763] = 32'h00000000,
        RAM[5764] = 32'h00000000,
        RAM[5765] = 32'h00000000,
        RAM[5766] = 32'h00000000,
        RAM[5767] = 32'h00000000,
        RAM[5768] = 32'h00000000,
        RAM[5769] = 32'h00000000,
        RAM[5770] = 32'h00000000,
        RAM[5771] = 32'h00000000,
        RAM[5772] = 32'h00000000,
        RAM[5773] = 32'h00000000,
        RAM[5774] = 32'h00000000,
        RAM[5775] = 32'h00000000,
        RAM[5776] = 32'h00000000,
        RAM[5777] = 32'h00000000,
        RAM[5778] = 32'h00000000,
        RAM[5779] = 32'h00000000,
        RAM[5780] = 32'h00000000,
        RAM[5781] = 32'h00000000,
        RAM[5782] = 32'h00000000,
        RAM[5783] = 32'h00000000,
        RAM[5784] = 32'h00000000,
        RAM[5785] = 32'h00000000,
        RAM[5786] = 32'h00000000,
        RAM[5787] = 32'h00000000,
        RAM[5788] = 32'h00000000,
        RAM[5789] = 32'h00000000,
        RAM[5790] = 32'h00000000,
        RAM[5791] = 32'h00000000,
        RAM[5792] = 32'h00000000,
        RAM[5793] = 32'h00000000,
        RAM[5794] = 32'h00000000,
        RAM[5795] = 32'h00000000,
        RAM[5796] = 32'h00000000,
        RAM[5797] = 32'h00000000,
        RAM[5798] = 32'h00000000,
        RAM[5799] = 32'h00000000,
        RAM[5800] = 32'h00000000,
        RAM[5801] = 32'h00000000,
        RAM[5802] = 32'h00000000,
        RAM[5803] = 32'h00000000,
        RAM[5804] = 32'h00000000,
        RAM[5805] = 32'h00000000,
        RAM[5806] = 32'h00000000,
        RAM[5807] = 32'h00000000,
        RAM[5808] = 32'h00000000,
        RAM[5809] = 32'h00000000,
        RAM[5810] = 32'h00000000,
        RAM[5811] = 32'h00000000,
        RAM[5812] = 32'h00000000,
        RAM[5813] = 32'h00000000,
        RAM[5814] = 32'h00000000,
        RAM[5815] = 32'h00000000,
        RAM[5816] = 32'h00000000,
        RAM[5817] = 32'h00000000,
        RAM[5818] = 32'h00000000,
        RAM[5819] = 32'h00000000,
        RAM[5820] = 32'h00000000,
        RAM[5821] = 32'h00000000,
        RAM[5822] = 32'h00000000,
        RAM[5823] = 32'h00000000,
        RAM[5824] = 32'h00000000,
        RAM[5825] = 32'h00000000,
        RAM[5826] = 32'h00000000,
        RAM[5827] = 32'h00000000,
        RAM[5828] = 32'h00000000,
        RAM[5829] = 32'h00000000,
        RAM[5830] = 32'h00000000,
        RAM[5831] = 32'h00000000,
        RAM[5832] = 32'h00000000,
        RAM[5833] = 32'h00000000,
        RAM[5834] = 32'h00000000,
        RAM[5835] = 32'h00000000,
        RAM[5836] = 32'h00000000,
        RAM[5837] = 32'h00000000,
        RAM[5838] = 32'h00000000,
        RAM[5839] = 32'h00000000,
        RAM[5840] = 32'h00000000,
        RAM[5841] = 32'h00000000,
        RAM[5842] = 32'h00000000,
        RAM[5843] = 32'h00000000,
        RAM[5844] = 32'h00000000,
        RAM[5845] = 32'h00000000,
        RAM[5846] = 32'h00000000,
        RAM[5847] = 32'h00000000,
        RAM[5848] = 32'h00000000,
        RAM[5849] = 32'h00000000,
        RAM[5850] = 32'h00000000,
        RAM[5851] = 32'h00000000,
        RAM[5852] = 32'h00000000,
        RAM[5853] = 32'h00000000,
        RAM[5854] = 32'h00000000,
        RAM[5855] = 32'h00000000,
        RAM[5856] = 32'h00000000,
        RAM[5857] = 32'h00000000,
        RAM[5858] = 32'h00000000,
        RAM[5859] = 32'h00000000,
        RAM[5860] = 32'h00000000,
        RAM[5861] = 32'h00000000,
        RAM[5862] = 32'h00000000,
        RAM[5863] = 32'h00000000,
        RAM[5864] = 32'h00000000,
        RAM[5865] = 32'h00000000,
        RAM[5866] = 32'h00000000,
        RAM[5867] = 32'h00000000,
        RAM[5868] = 32'h00000000,
        RAM[5869] = 32'h00000000,
        RAM[5870] = 32'h00000000,
        RAM[5871] = 32'h00000000,
        RAM[5872] = 32'h00000000,
        RAM[5873] = 32'h00000000,
        RAM[5874] = 32'h00000000,
        RAM[5875] = 32'h00000000,
        RAM[5876] = 32'h00000000,
        RAM[5877] = 32'h00000000,
        RAM[5878] = 32'h00000000,
        RAM[5879] = 32'h00000000,
        RAM[5880] = 32'h00000000,
        RAM[5881] = 32'h00000000,
        RAM[5882] = 32'h00000000,
        RAM[5883] = 32'h00000000,
        RAM[5884] = 32'h00000000,
        RAM[5885] = 32'h00000000,
        RAM[5886] = 32'h00000000,
        RAM[5887] = 32'h00000000,
        RAM[5888] = 32'h00000000,
        RAM[5889] = 32'h00000000,
        RAM[5890] = 32'h00000000,
        RAM[5891] = 32'h00000000,
        RAM[5892] = 32'h00000000,
        RAM[5893] = 32'h00000000,
        RAM[5894] = 32'h00000000,
        RAM[5895] = 32'h00000000,
        RAM[5896] = 32'h00000000,
        RAM[5897] = 32'h00000000,
        RAM[5898] = 32'h00000000,
        RAM[5899] = 32'h00000000,
        RAM[5900] = 32'h00000000,
        RAM[5901] = 32'h00000000,
        RAM[5902] = 32'h00000000,
        RAM[5903] = 32'h00000000,
        RAM[5904] = 32'h00000000,
        RAM[5905] = 32'h00000000,
        RAM[5906] = 32'h00000000,
        RAM[5907] = 32'h00000000,
        RAM[5908] = 32'h00000000,
        RAM[5909] = 32'h00000000,
        RAM[5910] = 32'h00000000,
        RAM[5911] = 32'h00000000,
        RAM[5912] = 32'h00000000,
        RAM[5913] = 32'h00000000,
        RAM[5914] = 32'h00000000,
        RAM[5915] = 32'h00000000,
        RAM[5916] = 32'h00000000,
        RAM[5917] = 32'h00000000,
        RAM[5918] = 32'h00000000,
        RAM[5919] = 32'h00000000,
        RAM[5920] = 32'h00000000,
        RAM[5921] = 32'h00000000,
        RAM[5922] = 32'h00000000,
        RAM[5923] = 32'h00000000,
        RAM[5924] = 32'h00000000,
        RAM[5925] = 32'h00000000,
        RAM[5926] = 32'h00000000,
        RAM[5927] = 32'h00000000,
        RAM[5928] = 32'h00000000,
        RAM[5929] = 32'h00000000,
        RAM[5930] = 32'h00000000,
        RAM[5931] = 32'h00000000,
        RAM[5932] = 32'h00000000,
        RAM[5933] = 32'h00000000,
        RAM[5934] = 32'h00000000,
        RAM[5935] = 32'h00000000,
        RAM[5936] = 32'h00000000,
        RAM[5937] = 32'h00000000,
        RAM[5938] = 32'h00000000,
        RAM[5939] = 32'h00000000,
        RAM[5940] = 32'h00000000,
        RAM[5941] = 32'h00000000,
        RAM[5942] = 32'h00000000,
        RAM[5943] = 32'h00000000,
        RAM[5944] = 32'h00000000,
        RAM[5945] = 32'h00000000,
        RAM[5946] = 32'h00000000,
        RAM[5947] = 32'h00000000,
        RAM[5948] = 32'h00000000,
        RAM[5949] = 32'h00000000,
        RAM[5950] = 32'h00000000,
        RAM[5951] = 32'h00000000,
        RAM[5952] = 32'h00000000,
        RAM[5953] = 32'h00000000,
        RAM[5954] = 32'h00000000,
        RAM[5955] = 32'h00000000,
        RAM[5956] = 32'h00000000,
        RAM[5957] = 32'h00000000,
        RAM[5958] = 32'h00000000,
        RAM[5959] = 32'h00000000,
        RAM[5960] = 32'h00000000,
        RAM[5961] = 32'h00000000,
        RAM[5962] = 32'h00000000,
        RAM[5963] = 32'h00000000,
        RAM[5964] = 32'h00000000,
        RAM[5965] = 32'h00000000,
        RAM[5966] = 32'h00000000,
        RAM[5967] = 32'h00000000,
        RAM[5968] = 32'h00000000,
        RAM[5969] = 32'h00000000,
        RAM[5970] = 32'h00000000,
        RAM[5971] = 32'h00000000,
        RAM[5972] = 32'h00000000,
        RAM[5973] = 32'h00000000,
        RAM[5974] = 32'h00000000,
        RAM[5975] = 32'h00000000,
        RAM[5976] = 32'h00000000,
        RAM[5977] = 32'h00000000,
        RAM[5978] = 32'h00000000,
        RAM[5979] = 32'h00000000,
        RAM[5980] = 32'h00000000,
        RAM[5981] = 32'h00000000,
        RAM[5982] = 32'h00000000,
        RAM[5983] = 32'h00000000,
        RAM[5984] = 32'h00000000,
        RAM[5985] = 32'h00000000,
        RAM[5986] = 32'h00000000,
        RAM[5987] = 32'h00000000,
        RAM[5988] = 32'h00000000,
        RAM[5989] = 32'h00000000,
        RAM[5990] = 32'h00000000,
        RAM[5991] = 32'h00000000,
        RAM[5992] = 32'h00000000,
        RAM[5993] = 32'h00000000,
        RAM[5994] = 32'h00000000,
        RAM[5995] = 32'h00000000,
        RAM[5996] = 32'h00000000,
        RAM[5997] = 32'h00000000,
        RAM[5998] = 32'h00000000,
        RAM[5999] = 32'h00000000,
        RAM[6000] = 32'h00000000,
        RAM[6001] = 32'h00000000,
        RAM[6002] = 32'h00000000,
        RAM[6003] = 32'h00000000,
        RAM[6004] = 32'h00000000,
        RAM[6005] = 32'h00000000,
        RAM[6006] = 32'h00000000,
        RAM[6007] = 32'h00000000,
        RAM[6008] = 32'h00000000,
        RAM[6009] = 32'h00000000,
        RAM[6010] = 32'h00000000,
        RAM[6011] = 32'h00000000,
        RAM[6012] = 32'h00000000,
        RAM[6013] = 32'h00000000,
        RAM[6014] = 32'h00000000,
        RAM[6015] = 32'h00000000,
        RAM[6016] = 32'h00000000,
        RAM[6017] = 32'h00000000,
        RAM[6018] = 32'h00000000,
        RAM[6019] = 32'h00000000,
        RAM[6020] = 32'h00000000,
        RAM[6021] = 32'h00000000,
        RAM[6022] = 32'h00000000,
        RAM[6023] = 32'h00000000,
        RAM[6024] = 32'h00000000,
        RAM[6025] = 32'h00000000,
        RAM[6026] = 32'h00000000,
        RAM[6027] = 32'h00000000,
        RAM[6028] = 32'h00000000,
        RAM[6029] = 32'h00000000,
        RAM[6030] = 32'h00000000,
        RAM[6031] = 32'h00000000,
        RAM[6032] = 32'h00000000,
        RAM[6033] = 32'h00000000,
        RAM[6034] = 32'h00000000,
        RAM[6035] = 32'h00000000,
        RAM[6036] = 32'h00000000,
        RAM[6037] = 32'h00000000,
        RAM[6038] = 32'h00000000,
        RAM[6039] = 32'h00000000,
        RAM[6040] = 32'h00000000,
        RAM[6041] = 32'h00000000,
        RAM[6042] = 32'h00000000,
        RAM[6043] = 32'h00000000,
        RAM[6044] = 32'h00000000,
        RAM[6045] = 32'h00000000,
        RAM[6046] = 32'h00000000,
        RAM[6047] = 32'h00000000,
        RAM[6048] = 32'h00000000,
        RAM[6049] = 32'h00000000,
        RAM[6050] = 32'h00000000,
        RAM[6051] = 32'h00000000,
        RAM[6052] = 32'h00000000,
        RAM[6053] = 32'h00000000,
        RAM[6054] = 32'h00000000,
        RAM[6055] = 32'h00000000,
        RAM[6056] = 32'h00000000,
        RAM[6057] = 32'h00000000,
        RAM[6058] = 32'h00000000,
        RAM[6059] = 32'h00000000,
        RAM[6060] = 32'h00000000,
        RAM[6061] = 32'h00000000,
        RAM[6062] = 32'h00000000,
        RAM[6063] = 32'h00000000,
        RAM[6064] = 32'h00000000,
        RAM[6065] = 32'h00000000,
        RAM[6066] = 32'h00000000,
        RAM[6067] = 32'h00000000,
        RAM[6068] = 32'h00000000,
        RAM[6069] = 32'h00000000,
        RAM[6070] = 32'h00000000,
        RAM[6071] = 32'h00000000,
        RAM[6072] = 32'h00000000,
        RAM[6073] = 32'h00000000,
        RAM[6074] = 32'h00000000,
        RAM[6075] = 32'h00000000,
        RAM[6076] = 32'h00000000,
        RAM[6077] = 32'h00000000,
        RAM[6078] = 32'h00000000,
        RAM[6079] = 32'h00000000,
        RAM[6080] = 32'h00000000,
        RAM[6081] = 32'h00000000,
        RAM[6082] = 32'h00000000,
        RAM[6083] = 32'h00000000,
        RAM[6084] = 32'h00000000,
        RAM[6085] = 32'h00000000,
        RAM[6086] = 32'h00000000,
        RAM[6087] = 32'h00000000,
        RAM[6088] = 32'h00000000,
        RAM[6089] = 32'h00000000,
        RAM[6090] = 32'h00000000,
        RAM[6091] = 32'h00000000,
        RAM[6092] = 32'h00000000,
        RAM[6093] = 32'h00000000,
        RAM[6094] = 32'h00000000,
        RAM[6095] = 32'h00000000,
        RAM[6096] = 32'h00000000,
        RAM[6097] = 32'h00000000,
        RAM[6098] = 32'h00000000,
        RAM[6099] = 32'h00000000,
        RAM[6100] = 32'h00000000,
        RAM[6101] = 32'h00000000,
        RAM[6102] = 32'h00000000,
        RAM[6103] = 32'h00000000,
        RAM[6104] = 32'h00000000,
        RAM[6105] = 32'h00000000,
        RAM[6106] = 32'h00000000,
        RAM[6107] = 32'h00000000,
        RAM[6108] = 32'h00000000,
        RAM[6109] = 32'h00000000,
        RAM[6110] = 32'h00000000,
        RAM[6111] = 32'h00000000,
        RAM[6112] = 32'h00000000,
        RAM[6113] = 32'h00000000,
        RAM[6114] = 32'h00000000,
        RAM[6115] = 32'h00000000,
        RAM[6116] = 32'h00000000,
        RAM[6117] = 32'h00000000,
        RAM[6118] = 32'h00000000,
        RAM[6119] = 32'h00000000,
        RAM[6120] = 32'h00000000,
        RAM[6121] = 32'h00000000,
        RAM[6122] = 32'h00000000,
        RAM[6123] = 32'h00000000,
        RAM[6124] = 32'h00000000,
        RAM[6125] = 32'h00000000,
        RAM[6126] = 32'h00000000,
        RAM[6127] = 32'h00000000,
        RAM[6128] = 32'h00000000,
        RAM[6129] = 32'h00000000,
        RAM[6130] = 32'h00000000,
        RAM[6131] = 32'h00000000,
        RAM[6132] = 32'h00000000,
        RAM[6133] = 32'h00000000,
        RAM[6134] = 32'h00000000,
        RAM[6135] = 32'h00000000,
        RAM[6136] = 32'h00000000,
        RAM[6137] = 32'h00000000,
        RAM[6138] = 32'h00000000,
        RAM[6139] = 32'h00000000,
        RAM[6140] = 32'h00000000,
        RAM[6141] = 32'h00000000,
        RAM[6142] = 32'h00000000,
        RAM[6143] = 32'h00000000,
        RAM[6144] = 32'h00000000,
        RAM[6145] = 32'h00000000,
        RAM[6146] = 32'h00000000,
        RAM[6147] = 32'h00000000,
        RAM[6148] = 32'h00000000,
        RAM[6149] = 32'h00000000,
        RAM[6150] = 32'h00000000,
        RAM[6151] = 32'h00000000,
        RAM[6152] = 32'h00000000,
        RAM[6153] = 32'h00000000,
        RAM[6154] = 32'h00000000,
        RAM[6155] = 32'h00000000,
        RAM[6156] = 32'h00000000,
        RAM[6157] = 32'h00000000,
        RAM[6158] = 32'h00000000,
        RAM[6159] = 32'h00000000,
        RAM[6160] = 32'h00000000,
        RAM[6161] = 32'h00000000,
        RAM[6162] = 32'h00000000,
        RAM[6163] = 32'h00000000,
        RAM[6164] = 32'h00000000,
        RAM[6165] = 32'h00000000,
        RAM[6166] = 32'h00000000,
        RAM[6167] = 32'h00000000,
        RAM[6168] = 32'h00000000,
        RAM[6169] = 32'h00000000,
        RAM[6170] = 32'h00000000,
        RAM[6171] = 32'h00000000,
        RAM[6172] = 32'h00000000,
        RAM[6173] = 32'h00000000,
        RAM[6174] = 32'h00000000,
        RAM[6175] = 32'h00000000,
        RAM[6176] = 32'h00000000,
        RAM[6177] = 32'h00000000,
        RAM[6178] = 32'h00000000,
        RAM[6179] = 32'h00000000,
        RAM[6180] = 32'h00000000,
        RAM[6181] = 32'h00000000,
        RAM[6182] = 32'h00000000,
        RAM[6183] = 32'h00000000,
        RAM[6184] = 32'h00000000,
        RAM[6185] = 32'h00000000,
        RAM[6186] = 32'h00000000,
        RAM[6187] = 32'h00000000,
        RAM[6188] = 32'h00000000,
        RAM[6189] = 32'h00000000,
        RAM[6190] = 32'h00000000,
        RAM[6191] = 32'h00000000,
        RAM[6192] = 32'h00000000,
        RAM[6193] = 32'h00000000,
        RAM[6194] = 32'h00000000,
        RAM[6195] = 32'h00000000,
        RAM[6196] = 32'h00000000,
        RAM[6197] = 32'h00000000,
        RAM[6198] = 32'h00000000,
        RAM[6199] = 32'h00000000,
        RAM[6200] = 32'h00000000,
        RAM[6201] = 32'h00000000,
        RAM[6202] = 32'h00000000,
        RAM[6203] = 32'h00000000,
        RAM[6204] = 32'h00000000,
        RAM[6205] = 32'h00000000,
        RAM[6206] = 32'h00000000,
        RAM[6207] = 32'h00000000,
        RAM[6208] = 32'h00000000,
        RAM[6209] = 32'h00000000,
        RAM[6210] = 32'h00000000,
        RAM[6211] = 32'h00000000,
        RAM[6212] = 32'h00000000,
        RAM[6213] = 32'h00000000,
        RAM[6214] = 32'h00000000,
        RAM[6215] = 32'h00000000,
        RAM[6216] = 32'h00000000,
        RAM[6217] = 32'h00000000,
        RAM[6218] = 32'h00000000,
        RAM[6219] = 32'h00000000,
        RAM[6220] = 32'h00000000,
        RAM[6221] = 32'h00000000,
        RAM[6222] = 32'h00000000,
        RAM[6223] = 32'h00000000,
        RAM[6224] = 32'h00000000,
        RAM[6225] = 32'h00000000,
        RAM[6226] = 32'h00000000,
        RAM[6227] = 32'h00000000,
        RAM[6228] = 32'h00000000,
        RAM[6229] = 32'h00000000,
        RAM[6230] = 32'h00000000,
        RAM[6231] = 32'h00000000,
        RAM[6232] = 32'h00000000,
        RAM[6233] = 32'h00000000,
        RAM[6234] = 32'h00000000,
        RAM[6235] = 32'h00000000,
        RAM[6236] = 32'h00000000,
        RAM[6237] = 32'h00000000,
        RAM[6238] = 32'h00000000,
        RAM[6239] = 32'h00000000,
        RAM[6240] = 32'h00000000,
        RAM[6241] = 32'h00000000,
        RAM[6242] = 32'h00000000,
        RAM[6243] = 32'h00000000,
        RAM[6244] = 32'h00000000,
        RAM[6245] = 32'h00000000,
        RAM[6246] = 32'h00000000,
        RAM[6247] = 32'h00000000,
        RAM[6248] = 32'h00000000,
        RAM[6249] = 32'h00000000,
        RAM[6250] = 32'h00000000,
        RAM[6251] = 32'h00000000,
        RAM[6252] = 32'h00000000,
        RAM[6253] = 32'h00000000,
        RAM[6254] = 32'h00000000,
        RAM[6255] = 32'h00000000,
        RAM[6256] = 32'h00000000,
        RAM[6257] = 32'h00000000,
        RAM[6258] = 32'h00000000,
        RAM[6259] = 32'h00000000,
        RAM[6260] = 32'h00000000,
        RAM[6261] = 32'h00000000,
        RAM[6262] = 32'h00000000,
        RAM[6263] = 32'h00000000,
        RAM[6264] = 32'h00000000,
        RAM[6265] = 32'h00000000,
        RAM[6266] = 32'h00000000,
        RAM[6267] = 32'h00000000,
        RAM[6268] = 32'h00000000,
        RAM[6269] = 32'h00000000,
        RAM[6270] = 32'h00000000,
        RAM[6271] = 32'h00000000,
        RAM[6272] = 32'h00000000,
        RAM[6273] = 32'h00000000,
        RAM[6274] = 32'h00000000,
        RAM[6275] = 32'h00000000,
        RAM[6276] = 32'h00000000,
        RAM[6277] = 32'h00000000,
        RAM[6278] = 32'h00000000,
        RAM[6279] = 32'h00000000,
        RAM[6280] = 32'h00000000,
        RAM[6281] = 32'h00000000,
        RAM[6282] = 32'h00000000,
        RAM[6283] = 32'h00000000,
        RAM[6284] = 32'h00000000,
        RAM[6285] = 32'h00000000,
        RAM[6286] = 32'h00000000,
        RAM[6287] = 32'h00000000,
        RAM[6288] = 32'h00000000,
        RAM[6289] = 32'h00000000,
        RAM[6290] = 32'h00000000,
        RAM[6291] = 32'h00000000,
        RAM[6292] = 32'h00000000,
        RAM[6293] = 32'h00000000,
        RAM[6294] = 32'h00000000,
        RAM[6295] = 32'h00000000,
        RAM[6296] = 32'h00000000,
        RAM[6297] = 32'h00000000,
        RAM[6298] = 32'h00000000,
        RAM[6299] = 32'h00000000,
        RAM[6300] = 32'h00000000,
        RAM[6301] = 32'h00000000,
        RAM[6302] = 32'h00000000,
        RAM[6303] = 32'h00000000,
        RAM[6304] = 32'h00000000,
        RAM[6305] = 32'h00000000,
        RAM[6306] = 32'h00000000,
        RAM[6307] = 32'h00000000,
        RAM[6308] = 32'h00000000,
        RAM[6309] = 32'h00000000,
        RAM[6310] = 32'h00000000,
        RAM[6311] = 32'h00000000,
        RAM[6312] = 32'h00000000,
        RAM[6313] = 32'h00000000,
        RAM[6314] = 32'h00000000,
        RAM[6315] = 32'h00000000,
        RAM[6316] = 32'h00000000,
        RAM[6317] = 32'h00000000,
        RAM[6318] = 32'h00000000,
        RAM[6319] = 32'h00000000,
        RAM[6320] = 32'h00000000,
        RAM[6321] = 32'h00000000,
        RAM[6322] = 32'h00000000,
        RAM[6323] = 32'h00000000,
        RAM[6324] = 32'h00000000,
        RAM[6325] = 32'h00000000,
        RAM[6326] = 32'h00000000,
        RAM[6327] = 32'h00000000,
        RAM[6328] = 32'h00000000,
        RAM[6329] = 32'h00000000,
        RAM[6330] = 32'h00000000,
        RAM[6331] = 32'h00000000,
        RAM[6332] = 32'h00000000,
        RAM[6333] = 32'h00000000,
        RAM[6334] = 32'h00000000,
        RAM[6335] = 32'h00000000,
        RAM[6336] = 32'h00000000,
        RAM[6337] = 32'h00000000,
        RAM[6338] = 32'h00000000,
        RAM[6339] = 32'h00000000,
        RAM[6340] = 32'h00000000,
        RAM[6341] = 32'h00000000,
        RAM[6342] = 32'h00000000,
        RAM[6343] = 32'h00000000,
        RAM[6344] = 32'h00000000,
        RAM[6345] = 32'h00000000,
        RAM[6346] = 32'h00000000,
        RAM[6347] = 32'h00000000,
        RAM[6348] = 32'h00000000,
        RAM[6349] = 32'h00000000,
        RAM[6350] = 32'h00000000,
        RAM[6351] = 32'h00000000,
        RAM[6352] = 32'h00000000,
        RAM[6353] = 32'h00000000,
        RAM[6354] = 32'h00000000,
        RAM[6355] = 32'h00000000,
        RAM[6356] = 32'h00000000,
        RAM[6357] = 32'h00000000,
        RAM[6358] = 32'h00000000,
        RAM[6359] = 32'h00000000,
        RAM[6360] = 32'h00000000,
        RAM[6361] = 32'h00000000,
        RAM[6362] = 32'h00000000,
        RAM[6363] = 32'h00000000,
        RAM[6364] = 32'h00000000,
        RAM[6365] = 32'h00000000,
        RAM[6366] = 32'h00000000,
        RAM[6367] = 32'h00000000,
        RAM[6368] = 32'h00000000,
        RAM[6369] = 32'h00000000,
        RAM[6370] = 32'h00000000,
        RAM[6371] = 32'h00000000,
        RAM[6372] = 32'h00000000,
        RAM[6373] = 32'h00000000,
        RAM[6374] = 32'h00000000,
        RAM[6375] = 32'h00000000,
        RAM[6376] = 32'h00000000,
        RAM[6377] = 32'h00000000,
        RAM[6378] = 32'h00000000,
        RAM[6379] = 32'h00000000,
        RAM[6380] = 32'h00000000,
        RAM[6381] = 32'h00000000,
        RAM[6382] = 32'h00000000,
        RAM[6383] = 32'h00000000,
        RAM[6384] = 32'h00000000,
        RAM[6385] = 32'h00000000,
        RAM[6386] = 32'h00000000,
        RAM[6387] = 32'h00000000,
        RAM[6388] = 32'h00000000,
        RAM[6389] = 32'h00000000,
        RAM[6390] = 32'h00000000,
        RAM[6391] = 32'h00000000,
        RAM[6392] = 32'h00000000,
        RAM[6393] = 32'h00000000,
        RAM[6394] = 32'h00000000,
        RAM[6395] = 32'h00000000,
        RAM[6396] = 32'h00000000,
        RAM[6397] = 32'h00000000,
        RAM[6398] = 32'h00000000,
        RAM[6399] = 32'h00000000,
        RAM[6400] = 32'h00000000,
        RAM[6401] = 32'h00000000,
        RAM[6402] = 32'h00000000,
        RAM[6403] = 32'h00000000,
        RAM[6404] = 32'h00000000,
        RAM[6405] = 32'h00000000,
        RAM[6406] = 32'h00000000,
        RAM[6407] = 32'h00000000,
        RAM[6408] = 32'h00000000,
        RAM[6409] = 32'h00000000,
        RAM[6410] = 32'h00000000,
        RAM[6411] = 32'h00000000,
        RAM[6412] = 32'h00000000,
        RAM[6413] = 32'h00000000,
        RAM[6414] = 32'h00000000,
        RAM[6415] = 32'h00000000,
        RAM[6416] = 32'h00000000,
        RAM[6417] = 32'h00000000,
        RAM[6418] = 32'h00000000,
        RAM[6419] = 32'h00000000,
        RAM[6420] = 32'h00000000,
        RAM[6421] = 32'h00000000,
        RAM[6422] = 32'h00000000,
        RAM[6423] = 32'h00000000,
        RAM[6424] = 32'h00000000,
        RAM[6425] = 32'h00000000,
        RAM[6426] = 32'h00000000,
        RAM[6427] = 32'h00000000,
        RAM[6428] = 32'h00000000,
        RAM[6429] = 32'h00000000,
        RAM[6430] = 32'h00000000,
        RAM[6431] = 32'h00000000,
        RAM[6432] = 32'h00000000,
        RAM[6433] = 32'h00000000,
        RAM[6434] = 32'h00000000,
        RAM[6435] = 32'h00000000,
        RAM[6436] = 32'h00000000,
        RAM[6437] = 32'h00000000,
        RAM[6438] = 32'h00000000,
        RAM[6439] = 32'h00000000,
        RAM[6440] = 32'h00000000,
        RAM[6441] = 32'h00000000,
        RAM[6442] = 32'h00000000,
        RAM[6443] = 32'h00000000,
        RAM[6444] = 32'h00000000,
        RAM[6445] = 32'h00000000,
        RAM[6446] = 32'h00000000,
        RAM[6447] = 32'h00000000,
        RAM[6448] = 32'h00000000,
        RAM[6449] = 32'h00000000,
        RAM[6450] = 32'h00000000,
        RAM[6451] = 32'h00000000,
        RAM[6452] = 32'h00000000,
        RAM[6453] = 32'h00000000,
        RAM[6454] = 32'h00000000,
        RAM[6455] = 32'h00000000,
        RAM[6456] = 32'h00000000,
        RAM[6457] = 32'h00000000,
        RAM[6458] = 32'h00000000,
        RAM[6459] = 32'h00000000,
        RAM[6460] = 32'h00000000,
        RAM[6461] = 32'h00000000,
        RAM[6462] = 32'h00000000,
        RAM[6463] = 32'h00000000,
        RAM[6464] = 32'h00000000,
        RAM[6465] = 32'h00000000,
        RAM[6466] = 32'h00000000,
        RAM[6467] = 32'h00000000,
        RAM[6468] = 32'h00000000,
        RAM[6469] = 32'h00000000,
        RAM[6470] = 32'h00000000,
        RAM[6471] = 32'h00000000,
        RAM[6472] = 32'h00000000,
        RAM[6473] = 32'h00000000,
        RAM[6474] = 32'h00000000,
        RAM[6475] = 32'h00000000,
        RAM[6476] = 32'h00000000,
        RAM[6477] = 32'h00000000,
        RAM[6478] = 32'h00000000,
        RAM[6479] = 32'h00000000,
        RAM[6480] = 32'h00000000,
        RAM[6481] = 32'h00000000,
        RAM[6482] = 32'h00000000,
        RAM[6483] = 32'h00000000,
        RAM[6484] = 32'h00000000,
        RAM[6485] = 32'h00000000,
        RAM[6486] = 32'h00000000,
        RAM[6487] = 32'h00000000,
        RAM[6488] = 32'h00000000,
        RAM[6489] = 32'h00000000,
        RAM[6490] = 32'h00000000,
        RAM[6491] = 32'h00000000,
        RAM[6492] = 32'h00000000,
        RAM[6493] = 32'h00000000,
        RAM[6494] = 32'h00000000,
        RAM[6495] = 32'h00000000,
        RAM[6496] = 32'h00000000,
        RAM[6497] = 32'h00000000,
        RAM[6498] = 32'h00000000,
        RAM[6499] = 32'h00000000,
        RAM[6500] = 32'h00000000,
        RAM[6501] = 32'h00000000,
        RAM[6502] = 32'h00000000,
        RAM[6503] = 32'h00000000,
        RAM[6504] = 32'h00000000,
        RAM[6505] = 32'h00000000,
        RAM[6506] = 32'h00000000,
        RAM[6507] = 32'h00000000,
        RAM[6508] = 32'h00000000,
        RAM[6509] = 32'h00000000,
        RAM[6510] = 32'h00000000,
        RAM[6511] = 32'h00000000,
        RAM[6512] = 32'h00000000,
        RAM[6513] = 32'h00000000,
        RAM[6514] = 32'h00000000,
        RAM[6515] = 32'h00000000,
        RAM[6516] = 32'h00000000,
        RAM[6517] = 32'h00000000,
        RAM[6518] = 32'h00000000,
        RAM[6519] = 32'h00000000,
        RAM[6520] = 32'h00000000,
        RAM[6521] = 32'h00000000,
        RAM[6522] = 32'h00000000,
        RAM[6523] = 32'h00000000,
        RAM[6524] = 32'h00000000,
        RAM[6525] = 32'h00000000,
        RAM[6526] = 32'h00000000,
        RAM[6527] = 32'h00000000,
        RAM[6528] = 32'h00000000,
        RAM[6529] = 32'h00000000,
        RAM[6530] = 32'h00000000,
        RAM[6531] = 32'h00000000,
        RAM[6532] = 32'h00000000,
        RAM[6533] = 32'h00000000,
        RAM[6534] = 32'h00000000,
        RAM[6535] = 32'h00000000,
        RAM[6536] = 32'h00000000,
        RAM[6537] = 32'h00000000,
        RAM[6538] = 32'h00000000,
        RAM[6539] = 32'h00000000,
        RAM[6540] = 32'h00000000,
        RAM[6541] = 32'h00000000,
        RAM[6542] = 32'h00000000,
        RAM[6543] = 32'h00000000,
        RAM[6544] = 32'h00000000,
        RAM[6545] = 32'h00000000,
        RAM[6546] = 32'h00000000,
        RAM[6547] = 32'h00000000,
        RAM[6548] = 32'h00000000,
        RAM[6549] = 32'h00000000,
        RAM[6550] = 32'h00000000,
        RAM[6551] = 32'h00000000,
        RAM[6552] = 32'h00000000,
        RAM[6553] = 32'h00000000,
        RAM[6554] = 32'h00000000,
        RAM[6555] = 32'h00000000,
        RAM[6556] = 32'h00000000,
        RAM[6557] = 32'h00000000,
        RAM[6558] = 32'h00000000,
        RAM[6559] = 32'h00000000,
        RAM[6560] = 32'h00000000,
        RAM[6561] = 32'h00000000,
        RAM[6562] = 32'h00000000,
        RAM[6563] = 32'h00000000,
        RAM[6564] = 32'h00000000,
        RAM[6565] = 32'h00000000,
        RAM[6566] = 32'h00000000,
        RAM[6567] = 32'h00000000,
        RAM[6568] = 32'h00000000,
        RAM[6569] = 32'h00000000,
        RAM[6570] = 32'h00000000,
        RAM[6571] = 32'h00000000,
        RAM[6572] = 32'h00000000,
        RAM[6573] = 32'h00000000,
        RAM[6574] = 32'h00000000,
        RAM[6575] = 32'h00000000,
        RAM[6576] = 32'h00000000,
        RAM[6577] = 32'h00000000,
        RAM[6578] = 32'h00000000,
        RAM[6579] = 32'h00000000,
        RAM[6580] = 32'h00000000,
        RAM[6581] = 32'h00000000,
        RAM[6582] = 32'h00000000,
        RAM[6583] = 32'h00000000,
        RAM[6584] = 32'h00000000,
        RAM[6585] = 32'h00000000,
        RAM[6586] = 32'h00000000,
        RAM[6587] = 32'h00000000,
        RAM[6588] = 32'h00000000,
        RAM[6589] = 32'h00000000,
        RAM[6590] = 32'h00000000,
        RAM[6591] = 32'h00000000,
        RAM[6592] = 32'h00000000,
        RAM[6593] = 32'h00000000,
        RAM[6594] = 32'h00000000,
        RAM[6595] = 32'h00000000,
        RAM[6596] = 32'h00000000,
        RAM[6597] = 32'h00000000,
        RAM[6598] = 32'h00000000,
        RAM[6599] = 32'h00000000,
        RAM[6600] = 32'h00000000,
        RAM[6601] = 32'h00000000,
        RAM[6602] = 32'h00000000,
        RAM[6603] = 32'h00000000,
        RAM[6604] = 32'h00000000,
        RAM[6605] = 32'h00000000,
        RAM[6606] = 32'h00000000,
        RAM[6607] = 32'h00000000,
        RAM[6608] = 32'h00000000,
        RAM[6609] = 32'h00000000,
        RAM[6610] = 32'h00000000,
        RAM[6611] = 32'h00000000,
        RAM[6612] = 32'h00000000,
        RAM[6613] = 32'h00000000,
        RAM[6614] = 32'h00000000,
        RAM[6615] = 32'h00000000,
        RAM[6616] = 32'h00000000,
        RAM[6617] = 32'h00000000,
        RAM[6618] = 32'h00000000,
        RAM[6619] = 32'h00000000,
        RAM[6620] = 32'h00000000,
        RAM[6621] = 32'h00000000,
        RAM[6622] = 32'h00000000,
        RAM[6623] = 32'h00000000,
        RAM[6624] = 32'h00000000,
        RAM[6625] = 32'h00000000,
        RAM[6626] = 32'h00000000,
        RAM[6627] = 32'h00000000,
        RAM[6628] = 32'h00000000,
        RAM[6629] = 32'h00000000,
        RAM[6630] = 32'h00000000,
        RAM[6631] = 32'h00000000,
        RAM[6632] = 32'h00000000,
        RAM[6633] = 32'h00000000,
        RAM[6634] = 32'h00000000,
        RAM[6635] = 32'h00000000,
        RAM[6636] = 32'h00000000,
        RAM[6637] = 32'h00000000,
        RAM[6638] = 32'h00000000,
        RAM[6639] = 32'h00000000,
        RAM[6640] = 32'h00000000,
        RAM[6641] = 32'h00000000,
        RAM[6642] = 32'h00000000,
        RAM[6643] = 32'h00000000,
        RAM[6644] = 32'h00000000,
        RAM[6645] = 32'h00000000,
        RAM[6646] = 32'h00000000,
        RAM[6647] = 32'h00000000,
        RAM[6648] = 32'h00000000,
        RAM[6649] = 32'h00000000,
        RAM[6650] = 32'h00000000,
        RAM[6651] = 32'h00000000,
        RAM[6652] = 32'h00000000,
        RAM[6653] = 32'h00000000,
        RAM[6654] = 32'h00000000,
        RAM[6655] = 32'h00000000,
        RAM[6656] = 32'h00000000,
        RAM[6657] = 32'h00000000,
        RAM[6658] = 32'h00000000,
        RAM[6659] = 32'h00000000,
        RAM[6660] = 32'h00000000,
        RAM[6661] = 32'h00000000,
        RAM[6662] = 32'h00000000,
        RAM[6663] = 32'h00000000,
        RAM[6664] = 32'h00000000,
        RAM[6665] = 32'h00000000,
        RAM[6666] = 32'h00000000,
        RAM[6667] = 32'h00000000,
        RAM[6668] = 32'h00000000,
        RAM[6669] = 32'h00000000,
        RAM[6670] = 32'h00000000,
        RAM[6671] = 32'h00000000,
        RAM[6672] = 32'h00000000,
        RAM[6673] = 32'h00000000,
        RAM[6674] = 32'h00000000,
        RAM[6675] = 32'h00000000,
        RAM[6676] = 32'h00000000,
        RAM[6677] = 32'h00000000,
        RAM[6678] = 32'h00000000,
        RAM[6679] = 32'h00000000,
        RAM[6680] = 32'h00000000,
        RAM[6681] = 32'h00000000,
        RAM[6682] = 32'h00000000,
        RAM[6683] = 32'h00000000,
        RAM[6684] = 32'h00000000,
        RAM[6685] = 32'h00000000,
        RAM[6686] = 32'h00000000,
        RAM[6687] = 32'h00000000,
        RAM[6688] = 32'h00000000,
        RAM[6689] = 32'h00000000,
        RAM[6690] = 32'h00000000,
        RAM[6691] = 32'h00000000,
        RAM[6692] = 32'h00000000,
        RAM[6693] = 32'h00000000,
        RAM[6694] = 32'h00000000,
        RAM[6695] = 32'h00000000,
        RAM[6696] = 32'h00000000,
        RAM[6697] = 32'h00000000,
        RAM[6698] = 32'h00000000,
        RAM[6699] = 32'h00000000,
        RAM[6700] = 32'h00000000,
        RAM[6701] = 32'h00000000,
        RAM[6702] = 32'h00000000,
        RAM[6703] = 32'h00000000,
        RAM[6704] = 32'h00000000,
        RAM[6705] = 32'h00000000,
        RAM[6706] = 32'h00000000,
        RAM[6707] = 32'h00000000,
        RAM[6708] = 32'h00000000,
        RAM[6709] = 32'h00000000,
        RAM[6710] = 32'h00000000,
        RAM[6711] = 32'h00000000,
        RAM[6712] = 32'h00000000,
        RAM[6713] = 32'h00000000,
        RAM[6714] = 32'h00000000,
        RAM[6715] = 32'h00000000,
        RAM[6716] = 32'h00000000,
        RAM[6717] = 32'h00000000,
        RAM[6718] = 32'h00000000,
        RAM[6719] = 32'h00000000,
        RAM[6720] = 32'h00000000,
        RAM[6721] = 32'h00000000,
        RAM[6722] = 32'h00000000,
        RAM[6723] = 32'h00000000,
        RAM[6724] = 32'h00000000,
        RAM[6725] = 32'h00000000,
        RAM[6726] = 32'h00000000,
        RAM[6727] = 32'h00000000,
        RAM[6728] = 32'h00000000,
        RAM[6729] = 32'h00000000,
        RAM[6730] = 32'h00000000,
        RAM[6731] = 32'h00000000,
        RAM[6732] = 32'h00000000,
        RAM[6733] = 32'h00000000,
        RAM[6734] = 32'h00000000,
        RAM[6735] = 32'h00000000,
        RAM[6736] = 32'h00000000,
        RAM[6737] = 32'h00000000,
        RAM[6738] = 32'h00000000,
        RAM[6739] = 32'h00000000,
        RAM[6740] = 32'h00000000,
        RAM[6741] = 32'h00000000,
        RAM[6742] = 32'h00000000,
        RAM[6743] = 32'h00000000,
        RAM[6744] = 32'h00000000,
        RAM[6745] = 32'h00000000,
        RAM[6746] = 32'h00000000,
        RAM[6747] = 32'h00000000,
        RAM[6748] = 32'h00000000,
        RAM[6749] = 32'h00000000,
        RAM[6750] = 32'h00000000,
        RAM[6751] = 32'h00000000,
        RAM[6752] = 32'h00000000,
        RAM[6753] = 32'h00000000,
        RAM[6754] = 32'h00000000,
        RAM[6755] = 32'h00000000,
        RAM[6756] = 32'h00000000,
        RAM[6757] = 32'h00000000,
        RAM[6758] = 32'h00000000,
        RAM[6759] = 32'h00000000,
        RAM[6760] = 32'h00000000,
        RAM[6761] = 32'h00000000,
        RAM[6762] = 32'h00000000,
        RAM[6763] = 32'h00000000,
        RAM[6764] = 32'h00000000,
        RAM[6765] = 32'h00000000,
        RAM[6766] = 32'h00000000,
        RAM[6767] = 32'h00000000,
        RAM[6768] = 32'h00000000,
        RAM[6769] = 32'h00000000,
        RAM[6770] = 32'h00000000,
        RAM[6771] = 32'h00000000,
        RAM[6772] = 32'h00000000,
        RAM[6773] = 32'h00000000,
        RAM[6774] = 32'h00000000,
        RAM[6775] = 32'h00000000,
        RAM[6776] = 32'h00000000,
        RAM[6777] = 32'h00000000,
        RAM[6778] = 32'h00000000,
        RAM[6779] = 32'h00000000,
        RAM[6780] = 32'h00000000,
        RAM[6781] = 32'h00000000,
        RAM[6782] = 32'h00000000,
        RAM[6783] = 32'h00000000,
        RAM[6784] = 32'h00000000,
        RAM[6785] = 32'h00000000,
        RAM[6786] = 32'h00000000,
        RAM[6787] = 32'h00000000,
        RAM[6788] = 32'h00000000,
        RAM[6789] = 32'h00000000,
        RAM[6790] = 32'h00000000,
        RAM[6791] = 32'h00000000,
        RAM[6792] = 32'h00000000,
        RAM[6793] = 32'h00000000,
        RAM[6794] = 32'h00000000,
        RAM[6795] = 32'h00000000,
        RAM[6796] = 32'h00000000,
        RAM[6797] = 32'h00000000,
        RAM[6798] = 32'h00000000,
        RAM[6799] = 32'h00000000,
        RAM[6800] = 32'h00000000,
        RAM[6801] = 32'h00000000,
        RAM[6802] = 32'h00000000,
        RAM[6803] = 32'h00000000,
        RAM[6804] = 32'h00000000,
        RAM[6805] = 32'h00000000,
        RAM[6806] = 32'h00000000,
        RAM[6807] = 32'h00000000,
        RAM[6808] = 32'h00000000,
        RAM[6809] = 32'h00000000,
        RAM[6810] = 32'h00000000,
        RAM[6811] = 32'h00000000,
        RAM[6812] = 32'h00000000,
        RAM[6813] = 32'h00000000,
        RAM[6814] = 32'h00000000,
        RAM[6815] = 32'h00000000,
        RAM[6816] = 32'h00000000,
        RAM[6817] = 32'h00000000,
        RAM[6818] = 32'h00000000,
        RAM[6819] = 32'h00000000,
        RAM[6820] = 32'h00000000,
        RAM[6821] = 32'h00000000,
        RAM[6822] = 32'h00000000,
        RAM[6823] = 32'h00000000,
        RAM[6824] = 32'h00000000,
        RAM[6825] = 32'h00000000,
        RAM[6826] = 32'h00000000,
        RAM[6827] = 32'h00000000,
        RAM[6828] = 32'h00000000,
        RAM[6829] = 32'h00000000,
        RAM[6830] = 32'h00000000,
        RAM[6831] = 32'h00000000,
        RAM[6832] = 32'h00000000,
        RAM[6833] = 32'h00000000,
        RAM[6834] = 32'h00000000,
        RAM[6835] = 32'h00000000,
        RAM[6836] = 32'h00000000,
        RAM[6837] = 32'h00000000,
        RAM[6838] = 32'h00000000,
        RAM[6839] = 32'h00000000,
        RAM[6840] = 32'h00000000,
        RAM[6841] = 32'h00000000,
        RAM[6842] = 32'h00000000,
        RAM[6843] = 32'h00000000,
        RAM[6844] = 32'h00000000,
        RAM[6845] = 32'h00000000,
        RAM[6846] = 32'h00000000,
        RAM[6847] = 32'h00000000,
        RAM[6848] = 32'h00000000,
        RAM[6849] = 32'h00000000,
        RAM[6850] = 32'h00000000,
        RAM[6851] = 32'h00000000,
        RAM[6852] = 32'h00000000,
        RAM[6853] = 32'h00000000,
        RAM[6854] = 32'h00000000,
        RAM[6855] = 32'h00000000,
        RAM[6856] = 32'h00000000,
        RAM[6857] = 32'h00000000,
        RAM[6858] = 32'h00000000,
        RAM[6859] = 32'h00000000,
        RAM[6860] = 32'h00000000,
        RAM[6861] = 32'h00000000,
        RAM[6862] = 32'h00000000,
        RAM[6863] = 32'h00000000,
        RAM[6864] = 32'h00000000,
        RAM[6865] = 32'h00000000,
        RAM[6866] = 32'h00000000,
        RAM[6867] = 32'h00000000,
        RAM[6868] = 32'h00000000,
        RAM[6869] = 32'h00000000,
        RAM[6870] = 32'h00000000,
        RAM[6871] = 32'h00000000,
        RAM[6872] = 32'h00000000,
        RAM[6873] = 32'h00000000,
        RAM[6874] = 32'h00000000,
        RAM[6875] = 32'h00000000,
        RAM[6876] = 32'h00000000,
        RAM[6877] = 32'h00000000,
        RAM[6878] = 32'h00000000,
        RAM[6879] = 32'h00000000,
        RAM[6880] = 32'h00000000,
        RAM[6881] = 32'h00000000,
        RAM[6882] = 32'h00000000,
        RAM[6883] = 32'h00000000,
        RAM[6884] = 32'h00000000,
        RAM[6885] = 32'h00000000,
        RAM[6886] = 32'h00000000,
        RAM[6887] = 32'h00000000,
        RAM[6888] = 32'h00000000,
        RAM[6889] = 32'h00000000,
        RAM[6890] = 32'h00000000,
        RAM[6891] = 32'h00000000,
        RAM[6892] = 32'h00000000,
        RAM[6893] = 32'h00000000,
        RAM[6894] = 32'h00000000,
        RAM[6895] = 32'h00000000,
        RAM[6896] = 32'h00000000,
        RAM[6897] = 32'h00000000,
        RAM[6898] = 32'h00000000,
        RAM[6899] = 32'h00000000,
        RAM[6900] = 32'h00000000,
        RAM[6901] = 32'h00000000,
        RAM[6902] = 32'h00000000,
        RAM[6903] = 32'h00000000,
        RAM[6904] = 32'h00000000,
        RAM[6905] = 32'h00000000,
        RAM[6906] = 32'h00000000,
        RAM[6907] = 32'h00000000,
        RAM[6908] = 32'h00000000,
        RAM[6909] = 32'h00000000,
        RAM[6910] = 32'h00000000,
        RAM[6911] = 32'h00000000,
        RAM[6912] = 32'h00000000,
        RAM[6913] = 32'h00000000,
        RAM[6914] = 32'h00000000,
        RAM[6915] = 32'h00000000,
        RAM[6916] = 32'h00000000,
        RAM[6917] = 32'h00000000,
        RAM[6918] = 32'h00000000,
        RAM[6919] = 32'h00000000,
        RAM[6920] = 32'h00000000,
        RAM[6921] = 32'h00000000,
        RAM[6922] = 32'h00000000,
        RAM[6923] = 32'h00000000,
        RAM[6924] = 32'h00000000,
        RAM[6925] = 32'h00000000,
        RAM[6926] = 32'h00000000,
        RAM[6927] = 32'h00000000,
        RAM[6928] = 32'h00000000,
        RAM[6929] = 32'h00000000,
        RAM[6930] = 32'h00000000,
        RAM[6931] = 32'h00000000,
        RAM[6932] = 32'h00000000,
        RAM[6933] = 32'h00000000,
        RAM[6934] = 32'h00000000,
        RAM[6935] = 32'h00000000,
        RAM[6936] = 32'h00000000,
        RAM[6937] = 32'h00000000,
        RAM[6938] = 32'h00000000,
        RAM[6939] = 32'h00000000,
        RAM[6940] = 32'h00000000,
        RAM[6941] = 32'h00000000,
        RAM[6942] = 32'h00000000,
        RAM[6943] = 32'h00000000,
        RAM[6944] = 32'h00000000,
        RAM[6945] = 32'h00000000,
        RAM[6946] = 32'h00000000,
        RAM[6947] = 32'h00000000,
        RAM[6948] = 32'h00000000,
        RAM[6949] = 32'h00000000,
        RAM[6950] = 32'h00000000,
        RAM[6951] = 32'h00000000,
        RAM[6952] = 32'h00000000,
        RAM[6953] = 32'h00000000,
        RAM[6954] = 32'h00000000,
        RAM[6955] = 32'h00000000,
        RAM[6956] = 32'h00000000,
        RAM[6957] = 32'h00000000,
        RAM[6958] = 32'h00000000,
        RAM[6959] = 32'h00000000,
        RAM[6960] = 32'h00000000,
        RAM[6961] = 32'h00000000,
        RAM[6962] = 32'h00000000,
        RAM[6963] = 32'h00000000,
        RAM[6964] = 32'h00000000,
        RAM[6965] = 32'h00000000,
        RAM[6966] = 32'h00000000,
        RAM[6967] = 32'h00000000,
        RAM[6968] = 32'h00000000,
        RAM[6969] = 32'h00000000,
        RAM[6970] = 32'h00000000,
        RAM[6971] = 32'h00000000,
        RAM[6972] = 32'h00000000,
        RAM[6973] = 32'h00000000,
        RAM[6974] = 32'h00000000,
        RAM[6975] = 32'h00000000,
        RAM[6976] = 32'h00000000,
        RAM[6977] = 32'h00000000,
        RAM[6978] = 32'h00000000,
        RAM[6979] = 32'h00000000,
        RAM[6980] = 32'h00000000,
        RAM[6981] = 32'h00000000,
        RAM[6982] = 32'h00000000,
        RAM[6983] = 32'h00000000,
        RAM[6984] = 32'h00000000,
        RAM[6985] = 32'h00000000,
        RAM[6986] = 32'h00000000,
        RAM[6987] = 32'h00000000,
        RAM[6988] = 32'h00000000,
        RAM[6989] = 32'h00000000,
        RAM[6990] = 32'h00000000,
        RAM[6991] = 32'h00000000,
        RAM[6992] = 32'h00000000,
        RAM[6993] = 32'h00000000,
        RAM[6994] = 32'h00000000,
        RAM[6995] = 32'h00000000,
        RAM[6996] = 32'h00000000,
        RAM[6997] = 32'h00000000,
        RAM[6998] = 32'h00000000,
        RAM[6999] = 32'h00000000,
        RAM[7000] = 32'h00000000,
        RAM[7001] = 32'h00000000,
        RAM[7002] = 32'h00000000,
        RAM[7003] = 32'h00000000,
        RAM[7004] = 32'h00000000,
        RAM[7005] = 32'h00000000,
        RAM[7006] = 32'h00000000,
        RAM[7007] = 32'h00000000,
        RAM[7008] = 32'h00000000,
        RAM[7009] = 32'h00000000,
        RAM[7010] = 32'h00000000,
        RAM[7011] = 32'h00000000,
        RAM[7012] = 32'h00000000,
        RAM[7013] = 32'h00000000,
        RAM[7014] = 32'h00000000,
        RAM[7015] = 32'h00000000,
        RAM[7016] = 32'h00000000,
        RAM[7017] = 32'h00000000,
        RAM[7018] = 32'h00000000,
        RAM[7019] = 32'h00000000,
        RAM[7020] = 32'h00000000,
        RAM[7021] = 32'h00000000,
        RAM[7022] = 32'h00000000,
        RAM[7023] = 32'h00000000,
        RAM[7024] = 32'h00000000,
        RAM[7025] = 32'h00000000,
        RAM[7026] = 32'h00000000,
        RAM[7027] = 32'h00000000,
        RAM[7028] = 32'h00000000,
        RAM[7029] = 32'h00000000,
        RAM[7030] = 32'h00000000,
        RAM[7031] = 32'h00000000,
        RAM[7032] = 32'h00000000,
        RAM[7033] = 32'h00000000,
        RAM[7034] = 32'h00000000,
        RAM[7035] = 32'h00000000,
        RAM[7036] = 32'h00000000,
        RAM[7037] = 32'h00000000,
        RAM[7038] = 32'h00000000,
        RAM[7039] = 32'h00000000,
        RAM[7040] = 32'h00000000,
        RAM[7041] = 32'h00000000,
        RAM[7042] = 32'h00000000,
        RAM[7043] = 32'h00000000,
        RAM[7044] = 32'h00000000,
        RAM[7045] = 32'h00000000,
        RAM[7046] = 32'h00000000,
        RAM[7047] = 32'h00000000,
        RAM[7048] = 32'h00000000,
        RAM[7049] = 32'h00000000,
        RAM[7050] = 32'h00000000,
        RAM[7051] = 32'h00000000,
        RAM[7052] = 32'h00000000,
        RAM[7053] = 32'h00000000,
        RAM[7054] = 32'h00000000,
        RAM[7055] = 32'h00000000,
        RAM[7056] = 32'h00000000,
        RAM[7057] = 32'h00000000,
        RAM[7058] = 32'h00000000,
        RAM[7059] = 32'h00000000,
        RAM[7060] = 32'h00000000,
        RAM[7061] = 32'h00000000,
        RAM[7062] = 32'h00000000,
        RAM[7063] = 32'h00000000,
        RAM[7064] = 32'h00000000,
        RAM[7065] = 32'h00000000,
        RAM[7066] = 32'h00000000,
        RAM[7067] = 32'h00000000,
        RAM[7068] = 32'h00000000,
        RAM[7069] = 32'h00000000,
        RAM[7070] = 32'h00000000,
        RAM[7071] = 32'h00000000,
        RAM[7072] = 32'h00000000,
        RAM[7073] = 32'h00000000,
        RAM[7074] = 32'h00000000,
        RAM[7075] = 32'h00000000,
        RAM[7076] = 32'h00000000,
        RAM[7077] = 32'h00000000,
        RAM[7078] = 32'h00000000,
        RAM[7079] = 32'h00000000,
        RAM[7080] = 32'h00000000,
        RAM[7081] = 32'h00000000,
        RAM[7082] = 32'h00000000,
        RAM[7083] = 32'h00000000,
        RAM[7084] = 32'h00000000,
        RAM[7085] = 32'h00000000,
        RAM[7086] = 32'h00000000,
        RAM[7087] = 32'h00000000,
        RAM[7088] = 32'h00000000,
        RAM[7089] = 32'h00000000,
        RAM[7090] = 32'h00000000,
        RAM[7091] = 32'h00000000,
        RAM[7092] = 32'h00000000,
        RAM[7093] = 32'h00000000,
        RAM[7094] = 32'h00000000,
        RAM[7095] = 32'h00000000,
        RAM[7096] = 32'h00000000,
        RAM[7097] = 32'h00000000,
        RAM[7098] = 32'h00000000,
        RAM[7099] = 32'h00000000,
        RAM[7100] = 32'h00000000,
        RAM[7101] = 32'h00000000,
        RAM[7102] = 32'h00000000,
        RAM[7103] = 32'h00000000,
        RAM[7104] = 32'h00000000,
        RAM[7105] = 32'h00000000,
        RAM[7106] = 32'h00000000,
        RAM[7107] = 32'h00000000,
        RAM[7108] = 32'h00000000,
        RAM[7109] = 32'h00000000,
        RAM[7110] = 32'h00000000,
        RAM[7111] = 32'h00000000,
        RAM[7112] = 32'h00000000,
        RAM[7113] = 32'h00000000,
        RAM[7114] = 32'h00000000,
        RAM[7115] = 32'h00000000,
        RAM[7116] = 32'h00000000,
        RAM[7117] = 32'h00000000,
        RAM[7118] = 32'h00000000,
        RAM[7119] = 32'h00000000,
        RAM[7120] = 32'h00000000,
        RAM[7121] = 32'h00000000,
        RAM[7122] = 32'h00000000,
        RAM[7123] = 32'h00000000,
        RAM[7124] = 32'h00000000,
        RAM[7125] = 32'h00000000,
        RAM[7126] = 32'h00000000,
        RAM[7127] = 32'h00000000,
        RAM[7128] = 32'h00000000,
        RAM[7129] = 32'h00000000,
        RAM[7130] = 32'h00000000,
        RAM[7131] = 32'h00000000,
        RAM[7132] = 32'h00000000,
        RAM[7133] = 32'h00000000,
        RAM[7134] = 32'h00000000,
        RAM[7135] = 32'h00000000,
        RAM[7136] = 32'h00000000,
        RAM[7137] = 32'h00000000,
        RAM[7138] = 32'h00000000,
        RAM[7139] = 32'h00000000,
        RAM[7140] = 32'h00000000,
        RAM[7141] = 32'h00000000,
        RAM[7142] = 32'h00000000,
        RAM[7143] = 32'h00000000,
        RAM[7144] = 32'h00000000,
        RAM[7145] = 32'h00000000,
        RAM[7146] = 32'h00000000,
        RAM[7147] = 32'h00000000,
        RAM[7148] = 32'h00000000,
        RAM[7149] = 32'h00000000,
        RAM[7150] = 32'h00000000,
        RAM[7151] = 32'h00000000,
        RAM[7152] = 32'h00000000,
        RAM[7153] = 32'h00000000,
        RAM[7154] = 32'h00000000,
        RAM[7155] = 32'h00000000,
        RAM[7156] = 32'h00000000,
        RAM[7157] = 32'h00000000,
        RAM[7158] = 32'h00000000,
        RAM[7159] = 32'h00000000,
        RAM[7160] = 32'h00000000,
        RAM[7161] = 32'h00000000,
        RAM[7162] = 32'h00000000,
        RAM[7163] = 32'h00000000,
        RAM[7164] = 32'h00000000,
        RAM[7165] = 32'h00000000,
        RAM[7166] = 32'h00000000,
        RAM[7167] = 32'h00000000,
        RAM[7168] = 32'h00000000,
        RAM[7169] = 32'h00000000,
        RAM[7170] = 32'h00000000,
        RAM[7171] = 32'h00000000,
        RAM[7172] = 32'h00000000,
        RAM[7173] = 32'h00000000,
        RAM[7174] = 32'h00000000,
        RAM[7175] = 32'h00000000,
        RAM[7176] = 32'h00000000,
        RAM[7177] = 32'h00000000,
        RAM[7178] = 32'h00000000,
        RAM[7179] = 32'h00000000,
        RAM[7180] = 32'h00000000,
        RAM[7181] = 32'h00000000,
        RAM[7182] = 32'h00000000,
        RAM[7183] = 32'h00000000,
        RAM[7184] = 32'h00000000,
        RAM[7185] = 32'h00000000,
        RAM[7186] = 32'h00000000,
        RAM[7187] = 32'h00000000,
        RAM[7188] = 32'h00000000,
        RAM[7189] = 32'h00000000,
        RAM[7190] = 32'h00000000,
        RAM[7191] = 32'h00000000,
        RAM[7192] = 32'h00000000,
        RAM[7193] = 32'h00000000,
        RAM[7194] = 32'h00000000,
        RAM[7195] = 32'h00000000,
        RAM[7196] = 32'h00000000,
        RAM[7197] = 32'h00000000,
        RAM[7198] = 32'h00000000,
        RAM[7199] = 32'h00000000,
        RAM[7200] = 32'h00000000,
        RAM[7201] = 32'h00000000,
        RAM[7202] = 32'h00000000,
        RAM[7203] = 32'h00000000,
        RAM[7204] = 32'h00000000,
        RAM[7205] = 32'h00000000,
        RAM[7206] = 32'h00000000,
        RAM[7207] = 32'h00000000,
        RAM[7208] = 32'h00000000,
        RAM[7209] = 32'h00000000,
        RAM[7210] = 32'h00000000,
        RAM[7211] = 32'h00000000,
        RAM[7212] = 32'h00000000,
        RAM[7213] = 32'h00000000,
        RAM[7214] = 32'h00000000,
        RAM[7215] = 32'h00000000,
        RAM[7216] = 32'h00000000,
        RAM[7217] = 32'h00000000,
        RAM[7218] = 32'h00000000,
        RAM[7219] = 32'h00000000,
        RAM[7220] = 32'h00000000,
        RAM[7221] = 32'h00000000,
        RAM[7222] = 32'h00000000,
        RAM[7223] = 32'h00000000,
        RAM[7224] = 32'h00000000,
        RAM[7225] = 32'h00000000,
        RAM[7226] = 32'h00000000,
        RAM[7227] = 32'h00000000,
        RAM[7228] = 32'h00000000,
        RAM[7229] = 32'h00000000,
        RAM[7230] = 32'h00000000,
        RAM[7231] = 32'h00000000,
        RAM[7232] = 32'h00000000,
        RAM[7233] = 32'h00000000,
        RAM[7234] = 32'h00000000,
        RAM[7235] = 32'h00000000,
        RAM[7236] = 32'h00000000,
        RAM[7237] = 32'h00000000,
        RAM[7238] = 32'h00000000,
        RAM[7239] = 32'h00000000,
        RAM[7240] = 32'h00000000,
        RAM[7241] = 32'h00000000,
        RAM[7242] = 32'h00000000,
        RAM[7243] = 32'h00000000,
        RAM[7244] = 32'h00000000,
        RAM[7245] = 32'h00000000,
        RAM[7246] = 32'h00000000,
        RAM[7247] = 32'h00000000,
        RAM[7248] = 32'h00000000,
        RAM[7249] = 32'h00000000,
        RAM[7250] = 32'h00000000,
        RAM[7251] = 32'h00000000,
        RAM[7252] = 32'h00000000,
        RAM[7253] = 32'h00000000,
        RAM[7254] = 32'h00000000,
        RAM[7255] = 32'h00000000,
        RAM[7256] = 32'h00000000,
        RAM[7257] = 32'h00000000,
        RAM[7258] = 32'h00000000,
        RAM[7259] = 32'h00000000,
        RAM[7260] = 32'h00000000,
        RAM[7261] = 32'h00000000,
        RAM[7262] = 32'h00000000,
        RAM[7263] = 32'h00000000,
        RAM[7264] = 32'h00000000,
        RAM[7265] = 32'h00000000,
        RAM[7266] = 32'h00000000,
        RAM[7267] = 32'h00000000,
        RAM[7268] = 32'h00000000,
        RAM[7269] = 32'h00000000,
        RAM[7270] = 32'h00000000,
        RAM[7271] = 32'h00000000,
        RAM[7272] = 32'h00000000,
        RAM[7273] = 32'h00000000,
        RAM[7274] = 32'h00000000,
        RAM[7275] = 32'h00000000,
        RAM[7276] = 32'h00000000,
        RAM[7277] = 32'h00000000,
        RAM[7278] = 32'h00000000,
        RAM[7279] = 32'h00000000,
        RAM[7280] = 32'h00000000,
        RAM[7281] = 32'h00000000,
        RAM[7282] = 32'h00000000,
        RAM[7283] = 32'h00000000,
        RAM[7284] = 32'h00000000,
        RAM[7285] = 32'h00000000,
        RAM[7286] = 32'h00000000,
        RAM[7287] = 32'h00000000,
        RAM[7288] = 32'h00000000,
        RAM[7289] = 32'h00000000,
        RAM[7290] = 32'h00000000,
        RAM[7291] = 32'h00000000,
        RAM[7292] = 32'h00000000,
        RAM[7293] = 32'h00000000,
        RAM[7294] = 32'h00000000,
        RAM[7295] = 32'h00000000,
        RAM[7296] = 32'h00000000,
        RAM[7297] = 32'h00000000,
        RAM[7298] = 32'h00000000,
        RAM[7299] = 32'h00000000,
        RAM[7300] = 32'h00000000,
        RAM[7301] = 32'h00000000,
        RAM[7302] = 32'h00000000,
        RAM[7303] = 32'h00000000,
        RAM[7304] = 32'h00000000,
        RAM[7305] = 32'h00000000,
        RAM[7306] = 32'h00000000,
        RAM[7307] = 32'h00000000,
        RAM[7308] = 32'h00000000,
        RAM[7309] = 32'h00000000,
        RAM[7310] = 32'h00000000,
        RAM[7311] = 32'h00000000,
        RAM[7312] = 32'h00000000,
        RAM[7313] = 32'h00000000,
        RAM[7314] = 32'h00000000,
        RAM[7315] = 32'h00000000,
        RAM[7316] = 32'h00000000,
        RAM[7317] = 32'h00000000,
        RAM[7318] = 32'h00000000,
        RAM[7319] = 32'h00000000,
        RAM[7320] = 32'h00000000,
        RAM[7321] = 32'h00000000,
        RAM[7322] = 32'h00000000,
        RAM[7323] = 32'h00000000,
        RAM[7324] = 32'h00000000,
        RAM[7325] = 32'h00000000,
        RAM[7326] = 32'h00000000,
        RAM[7327] = 32'h00000000,
        RAM[7328] = 32'h00000000,
        RAM[7329] = 32'h00000000,
        RAM[7330] = 32'h00000000,
        RAM[7331] = 32'h00000000,
        RAM[7332] = 32'h00000000,
        RAM[7333] = 32'h00000000,
        RAM[7334] = 32'h00000000,
        RAM[7335] = 32'h00000000,
        RAM[7336] = 32'h00000000,
        RAM[7337] = 32'h00000000,
        RAM[7338] = 32'h00000000,
        RAM[7339] = 32'h00000000,
        RAM[7340] = 32'h00000000,
        RAM[7341] = 32'h00000000,
        RAM[7342] = 32'h00000000,
        RAM[7343] = 32'h00000000,
        RAM[7344] = 32'h00000000,
        RAM[7345] = 32'h00000000,
        RAM[7346] = 32'h00000000,
        RAM[7347] = 32'h00000000,
        RAM[7348] = 32'h00000000,
        RAM[7349] = 32'h00000000,
        RAM[7350] = 32'h00000000,
        RAM[7351] = 32'h00000000,
        RAM[7352] = 32'h00000000,
        RAM[7353] = 32'h00000000,
        RAM[7354] = 32'h00000000,
        RAM[7355] = 32'h00000000,
        RAM[7356] = 32'h00000000,
        RAM[7357] = 32'h00000000,
        RAM[7358] = 32'h00000000,
        RAM[7359] = 32'h00000000,
        RAM[7360] = 32'h00000000,
        RAM[7361] = 32'h00000000,
        RAM[7362] = 32'h00000000,
        RAM[7363] = 32'h00000000,
        RAM[7364] = 32'h00000000,
        RAM[7365] = 32'h00000000,
        RAM[7366] = 32'h00000000,
        RAM[7367] = 32'h00000000,
        RAM[7368] = 32'h00000000,
        RAM[7369] = 32'h00000000,
        RAM[7370] = 32'h00000000,
        RAM[7371] = 32'h00000000,
        RAM[7372] = 32'h00000000,
        RAM[7373] = 32'h00000000,
        RAM[7374] = 32'h00000000,
        RAM[7375] = 32'h00000000,
        RAM[7376] = 32'h00000000,
        RAM[7377] = 32'h00000000,
        RAM[7378] = 32'h00000000,
        RAM[7379] = 32'h00000000,
        RAM[7380] = 32'h00000000,
        RAM[7381] = 32'h00000000,
        RAM[7382] = 32'h00000000,
        RAM[7383] = 32'h00000000,
        RAM[7384] = 32'h00000000,
        RAM[7385] = 32'h00000000,
        RAM[7386] = 32'h00000000,
        RAM[7387] = 32'h00000000,
        RAM[7388] = 32'h00000000,
        RAM[7389] = 32'h00000000,
        RAM[7390] = 32'h00000000,
        RAM[7391] = 32'h00000000,
        RAM[7392] = 32'h00000000,
        RAM[7393] = 32'h00000000,
        RAM[7394] = 32'h00000000,
        RAM[7395] = 32'h00000000,
        RAM[7396] = 32'h00000000,
        RAM[7397] = 32'h00000000,
        RAM[7398] = 32'h00000000,
        RAM[7399] = 32'h00000000,
        RAM[7400] = 32'h00000000,
        RAM[7401] = 32'h00000000,
        RAM[7402] = 32'h00000000,
        RAM[7403] = 32'h00000000,
        RAM[7404] = 32'h00000000,
        RAM[7405] = 32'h00000000,
        RAM[7406] = 32'h00000000,
        RAM[7407] = 32'h00000000,
        RAM[7408] = 32'h00000000,
        RAM[7409] = 32'h00000000,
        RAM[7410] = 32'h00000000,
        RAM[7411] = 32'h00000000,
        RAM[7412] = 32'h00000000,
        RAM[7413] = 32'h00000000,
        RAM[7414] = 32'h00000000,
        RAM[7415] = 32'h00000000,
        RAM[7416] = 32'h00000000,
        RAM[7417] = 32'h00000000,
        RAM[7418] = 32'h00000000,
        RAM[7419] = 32'h00000000,
        RAM[7420] = 32'h00000000,
        RAM[7421] = 32'h00000000,
        RAM[7422] = 32'h00000000,
        RAM[7423] = 32'h00000000,
        RAM[7424] = 32'h00000000,
        RAM[7425] = 32'h00000000,
        RAM[7426] = 32'h00000000,
        RAM[7427] = 32'h00000000,
        RAM[7428] = 32'h00000000,
        RAM[7429] = 32'h00000000,
        RAM[7430] = 32'h00000000,
        RAM[7431] = 32'h00000000,
        RAM[7432] = 32'h00000000,
        RAM[7433] = 32'h00000000,
        RAM[7434] = 32'h00000000,
        RAM[7435] = 32'h00000000,
        RAM[7436] = 32'h00000000,
        RAM[7437] = 32'h00000000,
        RAM[7438] = 32'h00000000,
        RAM[7439] = 32'h00000000,
        RAM[7440] = 32'h00000000,
        RAM[7441] = 32'h00000000,
        RAM[7442] = 32'h00000000,
        RAM[7443] = 32'h00000000,
        RAM[7444] = 32'h00000000,
        RAM[7445] = 32'h00000000,
        RAM[7446] = 32'h00000000,
        RAM[7447] = 32'h00000000,
        RAM[7448] = 32'h00000000,
        RAM[7449] = 32'h00000000,
        RAM[7450] = 32'h00000000,
        RAM[7451] = 32'h00000000,
        RAM[7452] = 32'h00000000,
        RAM[7453] = 32'h00000000,
        RAM[7454] = 32'h00000000,
        RAM[7455] = 32'h00000000,
        RAM[7456] = 32'h00000000,
        RAM[7457] = 32'h00000000,
        RAM[7458] = 32'h00000000,
        RAM[7459] = 32'h00000000,
        RAM[7460] = 32'h00000000,
        RAM[7461] = 32'h00000000,
        RAM[7462] = 32'h00000000,
        RAM[7463] = 32'h00000000,
        RAM[7464] = 32'h00000000,
        RAM[7465] = 32'h00000000,
        RAM[7466] = 32'h00000000,
        RAM[7467] = 32'h00000000,
        RAM[7468] = 32'h00000000,
        RAM[7469] = 32'h00000000,
        RAM[7470] = 32'h00000000,
        RAM[7471] = 32'h00000000,
        RAM[7472] = 32'h00000000,
        RAM[7473] = 32'h00000000,
        RAM[7474] = 32'h00000000,
        RAM[7475] = 32'h00000000,
        RAM[7476] = 32'h00000000,
        RAM[7477] = 32'h00000000,
        RAM[7478] = 32'h00000000,
        RAM[7479] = 32'h00000000,
        RAM[7480] = 32'h00000000,
        RAM[7481] = 32'h00000000,
        RAM[7482] = 32'h00000000,
        RAM[7483] = 32'h00000000,
        RAM[7484] = 32'h00000000,
        RAM[7485] = 32'h00000000,
        RAM[7486] = 32'h00000000,
        RAM[7487] = 32'h00000000,
        RAM[7488] = 32'h00000000,
        RAM[7489] = 32'h00000000,
        RAM[7490] = 32'h00000000,
        RAM[7491] = 32'h00000000,
        RAM[7492] = 32'h00000000,
        RAM[7493] = 32'h00000000,
        RAM[7494] = 32'h00000000,
        RAM[7495] = 32'h00000000,
        RAM[7496] = 32'h00000000,
        RAM[7497] = 32'h00000000,
        RAM[7498] = 32'h00000000,
        RAM[7499] = 32'h00000000,
        RAM[7500] = 32'h00000000,
        RAM[7501] = 32'h00000000,
        RAM[7502] = 32'h00000000,
        RAM[7503] = 32'h00000000,
        RAM[7504] = 32'h00000000,
        RAM[7505] = 32'h00000000,
        RAM[7506] = 32'h00000000,
        RAM[7507] = 32'h00000000,
        RAM[7508] = 32'h00000000,
        RAM[7509] = 32'h00000000,
        RAM[7510] = 32'h00000000,
        RAM[7511] = 32'h00000000,
        RAM[7512] = 32'h00000000,
        RAM[7513] = 32'h00000000,
        RAM[7514] = 32'h00000000,
        RAM[7515] = 32'h00000000,
        RAM[7516] = 32'h00000000,
        RAM[7517] = 32'h00000000,
        RAM[7518] = 32'h00000000,
        RAM[7519] = 32'h00000000,
        RAM[7520] = 32'h00000000,
        RAM[7521] = 32'h00000000,
        RAM[7522] = 32'h00000000,
        RAM[7523] = 32'h00000000,
        RAM[7524] = 32'h00000000,
        RAM[7525] = 32'h00000000,
        RAM[7526] = 32'h00000000,
        RAM[7527] = 32'h00000000,
        RAM[7528] = 32'h00000000,
        RAM[7529] = 32'h00000000,
        RAM[7530] = 32'h00000000,
        RAM[7531] = 32'h00000000,
        RAM[7532] = 32'h00000000,
        RAM[7533] = 32'h00000000,
        RAM[7534] = 32'h00000000,
        RAM[7535] = 32'h00000000,
        RAM[7536] = 32'h00000000,
        RAM[7537] = 32'h00000000,
        RAM[7538] = 32'h00000000,
        RAM[7539] = 32'h00000000,
        RAM[7540] = 32'h00000000,
        RAM[7541] = 32'h00000000,
        RAM[7542] = 32'h00000000,
        RAM[7543] = 32'h00000000,
        RAM[7544] = 32'h00000000,
        RAM[7545] = 32'h00000000,
        RAM[7546] = 32'h00000000,
        RAM[7547] = 32'h00000000,
        RAM[7548] = 32'h00000000,
        RAM[7549] = 32'h00000000,
        RAM[7550] = 32'h00000000,
        RAM[7551] = 32'h00000000,
        RAM[7552] = 32'h00000000,
        RAM[7553] = 32'h00000000,
        RAM[7554] = 32'h00000000,
        RAM[7555] = 32'h00000000,
        RAM[7556] = 32'h00000000,
        RAM[7557] = 32'h00000000,
        RAM[7558] = 32'h00000000,
        RAM[7559] = 32'h00000000,
        RAM[7560] = 32'h00000000,
        RAM[7561] = 32'h00000000,
        RAM[7562] = 32'h00000000,
        RAM[7563] = 32'h00000000,
        RAM[7564] = 32'h00000000,
        RAM[7565] = 32'h00000000,
        RAM[7566] = 32'h00000000,
        RAM[7567] = 32'h00000000,
        RAM[7568] = 32'h00000000,
        RAM[7569] = 32'h00000000,
        RAM[7570] = 32'h00000000,
        RAM[7571] = 32'h00000000,
        RAM[7572] = 32'h00000000,
        RAM[7573] = 32'h00000000,
        RAM[7574] = 32'h00000000,
        RAM[7575] = 32'h00000000,
        RAM[7576] = 32'h00000000,
        RAM[7577] = 32'h00000000,
        RAM[7578] = 32'h00000000,
        RAM[7579] = 32'h00000000,
        RAM[7580] = 32'h00000000,
        RAM[7581] = 32'h00000000,
        RAM[7582] = 32'h00000000,
        RAM[7583] = 32'h00000000,
        RAM[7584] = 32'h00000000,
        RAM[7585] = 32'h00000000,
        RAM[7586] = 32'h00000000,
        RAM[7587] = 32'h00000000,
        RAM[7588] = 32'h00000000,
        RAM[7589] = 32'h00000000,
        RAM[7590] = 32'h00000000,
        RAM[7591] = 32'h00000000,
        RAM[7592] = 32'h00000000,
        RAM[7593] = 32'h00000000,
        RAM[7594] = 32'h00000000,
        RAM[7595] = 32'h00000000,
        RAM[7596] = 32'h00000000,
        RAM[7597] = 32'h00000000,
        RAM[7598] = 32'h00000000,
        RAM[7599] = 32'h00000000,
        RAM[7600] = 32'h00000000,
        RAM[7601] = 32'h00000000,
        RAM[7602] = 32'h00000000,
        RAM[7603] = 32'h00000000,
        RAM[7604] = 32'h00000000,
        RAM[7605] = 32'h00000000,
        RAM[7606] = 32'h00000000,
        RAM[7607] = 32'h00000000,
        RAM[7608] = 32'h00000000,
        RAM[7609] = 32'h00000000,
        RAM[7610] = 32'h00000000,
        RAM[7611] = 32'h00000000,
        RAM[7612] = 32'h00000000,
        RAM[7613] = 32'h00000000,
        RAM[7614] = 32'h00000000,
        RAM[7615] = 32'h00000000,
        RAM[7616] = 32'h00000000,
        RAM[7617] = 32'h00000000,
        RAM[7618] = 32'h00000000,
        RAM[7619] = 32'h00000000,
        RAM[7620] = 32'h00000000,
        RAM[7621] = 32'h00000000,
        RAM[7622] = 32'h00000000,
        RAM[7623] = 32'h00000000,
        RAM[7624] = 32'h00000000,
        RAM[7625] = 32'h00000000,
        RAM[7626] = 32'h00000000,
        RAM[7627] = 32'h00000000,
        RAM[7628] = 32'h00000000,
        RAM[7629] = 32'h00000000,
        RAM[7630] = 32'h00000000,
        RAM[7631] = 32'h00000000,
        RAM[7632] = 32'h00000000,
        RAM[7633] = 32'h00000000,
        RAM[7634] = 32'h00000000,
        RAM[7635] = 32'h00000000,
        RAM[7636] = 32'h00000000,
        RAM[7637] = 32'h00000000,
        RAM[7638] = 32'h00000000,
        RAM[7639] = 32'h00000000,
        RAM[7640] = 32'h00000000,
        RAM[7641] = 32'h00000000,
        RAM[7642] = 32'h00000000,
        RAM[7643] = 32'h00000000,
        RAM[7644] = 32'h00000000,
        RAM[7645] = 32'h00000000,
        RAM[7646] = 32'h00000000,
        RAM[7647] = 32'h00000000,
        RAM[7648] = 32'h00000000,
        RAM[7649] = 32'h00000000,
        RAM[7650] = 32'h00000000,
        RAM[7651] = 32'h00000000,
        RAM[7652] = 32'h00000000,
        RAM[7653] = 32'h00000000,
        RAM[7654] = 32'h00000000,
        RAM[7655] = 32'h00000000,
        RAM[7656] = 32'h00000000,
        RAM[7657] = 32'h00000000,
        RAM[7658] = 32'h00000000,
        RAM[7659] = 32'h00000000,
        RAM[7660] = 32'h00000000,
        RAM[7661] = 32'h00000000,
        RAM[7662] = 32'h00000000,
        RAM[7663] = 32'h00000000,
        RAM[7664] = 32'h00000000,
        RAM[7665] = 32'h00000000,
        RAM[7666] = 32'h00000000,
        RAM[7667] = 32'h00000000,
        RAM[7668] = 32'h00000000,
        RAM[7669] = 32'h00000000,
        RAM[7670] = 32'h00000000,
        RAM[7671] = 32'h00000000,
        RAM[7672] = 32'h00000000,
        RAM[7673] = 32'h00000000,
        RAM[7674] = 32'h00000000,
        RAM[7675] = 32'h00000000,
        RAM[7676] = 32'h00000000,
        RAM[7677] = 32'h00000000,
        RAM[7678] = 32'h00000000,
        RAM[7679] = 32'h00000000,
        RAM[7680] = 32'h00000000,
        RAM[7681] = 32'h00000000,
        RAM[7682] = 32'h00000000,
        RAM[7683] = 32'h00000000,
        RAM[7684] = 32'h00000000,
        RAM[7685] = 32'h00000000,
        RAM[7686] = 32'h00000000,
        RAM[7687] = 32'h00000000,
        RAM[7688] = 32'h00000000,
        RAM[7689] = 32'h00000000,
        RAM[7690] = 32'h00000000,
        RAM[7691] = 32'h00000000,
        RAM[7692] = 32'h00000000,
        RAM[7693] = 32'h00000000,
        RAM[7694] = 32'h00000000,
        RAM[7695] = 32'h00000000,
        RAM[7696] = 32'h00000000,
        RAM[7697] = 32'h00000000,
        RAM[7698] = 32'h00000000,
        RAM[7699] = 32'h00000000,
        RAM[7700] = 32'h00000000,
        RAM[7701] = 32'h00000000,
        RAM[7702] = 32'h00000000,
        RAM[7703] = 32'h00000000,
        RAM[7704] = 32'h00000000,
        RAM[7705] = 32'h00000000,
        RAM[7706] = 32'h00000000,
        RAM[7707] = 32'h00000000,
        RAM[7708] = 32'h00000000,
        RAM[7709] = 32'h00000000,
        RAM[7710] = 32'h00000000,
        RAM[7711] = 32'h00000000,
        RAM[7712] = 32'h00000000,
        RAM[7713] = 32'h00000000,
        RAM[7714] = 32'h00000000,
        RAM[7715] = 32'h00000000,
        RAM[7716] = 32'h00000000,
        RAM[7717] = 32'h00000000,
        RAM[7718] = 32'h00000000,
        RAM[7719] = 32'h00000000,
        RAM[7720] = 32'h00000000,
        RAM[7721] = 32'h00000000,
        RAM[7722] = 32'h00000000,
        RAM[7723] = 32'h00000000,
        RAM[7724] = 32'h00000000,
        RAM[7725] = 32'h00000000,
        RAM[7726] = 32'h00000000,
        RAM[7727] = 32'h00000000,
        RAM[7728] = 32'h00000000,
        RAM[7729] = 32'h00000000,
        RAM[7730] = 32'h00000000,
        RAM[7731] = 32'h00000000,
        RAM[7732] = 32'h00000000,
        RAM[7733] = 32'h00000000,
        RAM[7734] = 32'h00000000,
        RAM[7735] = 32'h00000000,
        RAM[7736] = 32'h00000000,
        RAM[7737] = 32'h00000000,
        RAM[7738] = 32'h00000000,
        RAM[7739] = 32'h00000000,
        RAM[7740] = 32'h00000000,
        RAM[7741] = 32'h00000000,
        RAM[7742] = 32'h00000000,
        RAM[7743] = 32'h00000000,
        RAM[7744] = 32'h00000000,
        RAM[7745] = 32'h00000000,
        RAM[7746] = 32'h00000000,
        RAM[7747] = 32'h00000000,
        RAM[7748] = 32'h00000000,
        RAM[7749] = 32'h00000000,
        RAM[7750] = 32'h00000000,
        RAM[7751] = 32'h00000000,
        RAM[7752] = 32'h00000000,
        RAM[7753] = 32'h00000000,
        RAM[7754] = 32'h00000000,
        RAM[7755] = 32'h00000000,
        RAM[7756] = 32'h00000000,
        RAM[7757] = 32'h00000000,
        RAM[7758] = 32'h00000000,
        RAM[7759] = 32'h00000000,
        RAM[7760] = 32'h00000000,
        RAM[7761] = 32'h00000000,
        RAM[7762] = 32'h00000000,
        RAM[7763] = 32'h00000000,
        RAM[7764] = 32'h00000000,
        RAM[7765] = 32'h00000000,
        RAM[7766] = 32'h00000000,
        RAM[7767] = 32'h00000000,
        RAM[7768] = 32'h00000000,
        RAM[7769] = 32'h00000000,
        RAM[7770] = 32'h00000000,
        RAM[7771] = 32'h00000000,
        RAM[7772] = 32'h00000000,
        RAM[7773] = 32'h00000000,
        RAM[7774] = 32'h00000000,
        RAM[7775] = 32'h00000000,
        RAM[7776] = 32'h00000000,
        RAM[7777] = 32'h00000000,
        RAM[7778] = 32'h00000000,
        RAM[7779] = 32'h00000000,
        RAM[7780] = 32'h00000000,
        RAM[7781] = 32'h00000000,
        RAM[7782] = 32'h00000000,
        RAM[7783] = 32'h00000000,
        RAM[7784] = 32'h00000000,
        RAM[7785] = 32'h00000000,
        RAM[7786] = 32'h00000000,
        RAM[7787] = 32'h00000000,
        RAM[7788] = 32'h00000000,
        RAM[7789] = 32'h00000000,
        RAM[7790] = 32'h00000000,
        RAM[7791] = 32'h00000000,
        RAM[7792] = 32'h00000000,
        RAM[7793] = 32'h00000000,
        RAM[7794] = 32'h00000000,
        RAM[7795] = 32'h00000000,
        RAM[7796] = 32'h00000000,
        RAM[7797] = 32'h00000000,
        RAM[7798] = 32'h00000000,
        RAM[7799] = 32'h00000000,
        RAM[7800] = 32'h00000000,
        RAM[7801] = 32'h00000000,
        RAM[7802] = 32'h00000000,
        RAM[7803] = 32'h00000000,
        RAM[7804] = 32'h00000000,
        RAM[7805] = 32'h00000000,
        RAM[7806] = 32'h00000000,
        RAM[7807] = 32'h00000000,
        RAM[7808] = 32'h00000000,
        RAM[7809] = 32'h00000000,
        RAM[7810] = 32'h00000000,
        RAM[7811] = 32'h00000000,
        RAM[7812] = 32'h00000000,
        RAM[7813] = 32'h00000000,
        RAM[7814] = 32'h00000000,
        RAM[7815] = 32'h00000000,
        RAM[7816] = 32'h00000000,
        RAM[7817] = 32'h00000000,
        RAM[7818] = 32'h00000000,
        RAM[7819] = 32'h00000000,
        RAM[7820] = 32'h00000000,
        RAM[7821] = 32'h00000000,
        RAM[7822] = 32'h00000000,
        RAM[7823] = 32'h00000000,
        RAM[7824] = 32'h00000000,
        RAM[7825] = 32'h00000000,
        RAM[7826] = 32'h00000000,
        RAM[7827] = 32'h00000000,
        RAM[7828] = 32'h00000000,
        RAM[7829] = 32'h00000000,
        RAM[7830] = 32'h00000000,
        RAM[7831] = 32'h00000000,
        RAM[7832] = 32'h00000000,
        RAM[7833] = 32'h00000000,
        RAM[7834] = 32'h00000000,
        RAM[7835] = 32'h00000000,
        RAM[7836] = 32'h00000000,
        RAM[7837] = 32'h00000000,
        RAM[7838] = 32'h00000000,
        RAM[7839] = 32'h00000000,
        RAM[7840] = 32'h00000000,
        RAM[7841] = 32'h00000000,
        RAM[7842] = 32'h00000000,
        RAM[7843] = 32'h00000000,
        RAM[7844] = 32'h00000000,
        RAM[7845] = 32'h00000000,
        RAM[7846] = 32'h00000000,
        RAM[7847] = 32'h00000000,
        RAM[7848] = 32'h00000000,
        RAM[7849] = 32'h00000000,
        RAM[7850] = 32'h00000000,
        RAM[7851] = 32'h00000000,
        RAM[7852] = 32'h00000000,
        RAM[7853] = 32'h00000000,
        RAM[7854] = 32'h00000000,
        RAM[7855] = 32'h00000000,
        RAM[7856] = 32'h00000000,
        RAM[7857] = 32'h00000000,
        RAM[7858] = 32'h00000000,
        RAM[7859] = 32'h00000000,
        RAM[7860] = 32'h00000000,
        RAM[7861] = 32'h00000000,
        RAM[7862] = 32'h00000000,
        RAM[7863] = 32'h00000000,
        RAM[7864] = 32'h00000000,
        RAM[7865] = 32'h00000000,
        RAM[7866] = 32'h00000000,
        RAM[7867] = 32'h00000000,
        RAM[7868] = 32'h00000000,
        RAM[7869] = 32'h00000000,
        RAM[7870] = 32'h00000000,
        RAM[7871] = 32'h00000000,
        RAM[7872] = 32'h00000000,
        RAM[7873] = 32'h00000000,
        RAM[7874] = 32'h00000000,
        RAM[7875] = 32'h00000000,
        RAM[7876] = 32'h00000000,
        RAM[7877] = 32'h00000000,
        RAM[7878] = 32'h00000000,
        RAM[7879] = 32'h00000000,
        RAM[7880] = 32'h00000000,
        RAM[7881] = 32'h00000000,
        RAM[7882] = 32'h00000000,
        RAM[7883] = 32'h00000000,
        RAM[7884] = 32'h00000000,
        RAM[7885] = 32'h00000000,
        RAM[7886] = 32'h00000000,
        RAM[7887] = 32'h00000000,
        RAM[7888] = 32'h00000000,
        RAM[7889] = 32'h00000000,
        RAM[7890] = 32'h00000000,
        RAM[7891] = 32'h00000000,
        RAM[7892] = 32'h00000000,
        RAM[7893] = 32'h00000000,
        RAM[7894] = 32'h00000000,
        RAM[7895] = 32'h00000000,
        RAM[7896] = 32'h00000000,
        RAM[7897] = 32'h00000000,
        RAM[7898] = 32'h00000000,
        RAM[7899] = 32'h00000000,
        RAM[7900] = 32'h00000000,
        RAM[7901] = 32'h00000000,
        RAM[7902] = 32'h00000000,
        RAM[7903] = 32'h00000000,
        RAM[7904] = 32'h00000000,
        RAM[7905] = 32'h00000000,
        RAM[7906] = 32'h00000000,
        RAM[7907] = 32'h00000000,
        RAM[7908] = 32'h00000000,
        RAM[7909] = 32'h00000000,
        RAM[7910] = 32'h00000000,
        RAM[7911] = 32'h00000000,
        RAM[7912] = 32'h00000000,
        RAM[7913] = 32'h00000000,
        RAM[7914] = 32'h00000000,
        RAM[7915] = 32'h00000000,
        RAM[7916] = 32'h00000000,
        RAM[7917] = 32'h00000000,
        RAM[7918] = 32'h00000000,
        RAM[7919] = 32'h00000000,
        RAM[7920] = 32'h00000000,
        RAM[7921] = 32'h00000000,
        RAM[7922] = 32'h00000000,
        RAM[7923] = 32'h00000000,
        RAM[7924] = 32'h00000000,
        RAM[7925] = 32'h00000000,
        RAM[7926] = 32'h00000000,
        RAM[7927] = 32'h00000000,
        RAM[7928] = 32'h00000000,
        RAM[7929] = 32'h00000000,
        RAM[7930] = 32'h00000000,
        RAM[7931] = 32'h00000000,
        RAM[7932] = 32'h00000000,
        RAM[7933] = 32'h00000000,
        RAM[7934] = 32'h00000000,
        RAM[7935] = 32'h00000000,
        RAM[7936] = 32'h00000000,
        RAM[7937] = 32'h00000000,
        RAM[7938] = 32'h00000000,
        RAM[7939] = 32'h00000000,
        RAM[7940] = 32'h00000000,
        RAM[7941] = 32'h00000000,
        RAM[7942] = 32'h00000000,
        RAM[7943] = 32'h00000000,
        RAM[7944] = 32'h00000000,
        RAM[7945] = 32'h00000000,
        RAM[7946] = 32'h00000000,
        RAM[7947] = 32'h00000000,
        RAM[7948] = 32'h00000000,
        RAM[7949] = 32'h00000000,
        RAM[7950] = 32'h00000000,
        RAM[7951] = 32'h00000000,
        RAM[7952] = 32'h00000000,
        RAM[7953] = 32'h00000000,
        RAM[7954] = 32'h00000000,
        RAM[7955] = 32'h00000000,
        RAM[7956] = 32'h00000000,
        RAM[7957] = 32'h00000000,
        RAM[7958] = 32'h00000000,
        RAM[7959] = 32'h00000000,
        RAM[7960] = 32'h00000000,
        RAM[7961] = 32'h00000000,
        RAM[7962] = 32'h00000000,
        RAM[7963] = 32'h00000000,
        RAM[7964] = 32'h00000000,
        RAM[7965] = 32'h00000000,
        RAM[7966] = 32'h00000000,
        RAM[7967] = 32'h00000000,
        RAM[7968] = 32'h00000000,
        RAM[7969] = 32'h00000000,
        RAM[7970] = 32'h00000000,
        RAM[7971] = 32'h00000000,
        RAM[7972] = 32'h00000000,
        RAM[7973] = 32'h00000000,
        RAM[7974] = 32'h00000000,
        RAM[7975] = 32'h00000000,
        RAM[7976] = 32'h00000000,
        RAM[7977] = 32'h00000000,
        RAM[7978] = 32'h00000000,
        RAM[7979] = 32'h00000000,
        RAM[7980] = 32'h00000000,
        RAM[7981] = 32'h00000000,
        RAM[7982] = 32'h00000000,
        RAM[7983] = 32'h00000000,
        RAM[7984] = 32'h00000000,
        RAM[7985] = 32'h00000000,
        RAM[7986] = 32'h00000000,
        RAM[7987] = 32'h00000000,
        RAM[7988] = 32'h00000000,
        RAM[7989] = 32'h00000000,
        RAM[7990] = 32'h00000000,
        RAM[7991] = 32'h00000000,
        RAM[7992] = 32'h00000000,
        RAM[7993] = 32'h00000000,
        RAM[7994] = 32'h00000000,
        RAM[7995] = 32'h00000000,
        RAM[7996] = 32'h00000000,
        RAM[7997] = 32'h00000000,
        RAM[7998] = 32'h00000000,
        RAM[7999] = 32'h00000000,
        RAM[8000] = 32'h00000000,
        RAM[8001] = 32'h00000000,
        RAM[8002] = 32'h00000000,
        RAM[8003] = 32'h00000000,
        RAM[8004] = 32'h00000000,
        RAM[8005] = 32'h00000000,
        RAM[8006] = 32'h00000000,
        RAM[8007] = 32'h00000000,
        RAM[8008] = 32'h00000000,
        RAM[8009] = 32'h00000000,
        RAM[8010] = 32'h00000000,
        RAM[8011] = 32'h00000000,
        RAM[8012] = 32'h00000000,
        RAM[8013] = 32'h00000000,
        RAM[8014] = 32'h00000000,
        RAM[8015] = 32'h00000000,
        RAM[8016] = 32'h00000000,
        RAM[8017] = 32'h00000000,
        RAM[8018] = 32'h00000000,
        RAM[8019] = 32'h00000000,
        RAM[8020] = 32'h00000000,
        RAM[8021] = 32'h00000000,
        RAM[8022] = 32'h00000000,
        RAM[8023] = 32'h00000000,
        RAM[8024] = 32'h00000000,
        RAM[8025] = 32'h00000000,
        RAM[8026] = 32'h00000000,
        RAM[8027] = 32'h00000000,
        RAM[8028] = 32'h00000000,
        RAM[8029] = 32'h00000000,
        RAM[8030] = 32'h00000000,
        RAM[8031] = 32'h00000000,
        RAM[8032] = 32'h00000000,
        RAM[8033] = 32'h00000000,
        RAM[8034] = 32'h00000000,
        RAM[8035] = 32'h00000000,
        RAM[8036] = 32'h00000000,
        RAM[8037] = 32'h00000000,
        RAM[8038] = 32'h00000000,
        RAM[8039] = 32'h00000000,
        RAM[8040] = 32'h00000000,
        RAM[8041] = 32'h00000000,
        RAM[8042] = 32'h00000000,
        RAM[8043] = 32'h00000000,
        RAM[8044] = 32'h00000000,
        RAM[8045] = 32'h00000000,
        RAM[8046] = 32'h00000000,
        RAM[8047] = 32'h00000000,
        RAM[8048] = 32'h00000000,
        RAM[8049] = 32'h00000000,
        RAM[8050] = 32'h00000000,
        RAM[8051] = 32'h00000000,
        RAM[8052] = 32'h00000000,
        RAM[8053] = 32'h00000000,
        RAM[8054] = 32'h00000000,
        RAM[8055] = 32'h00000000,
        RAM[8056] = 32'h00000000,
        RAM[8057] = 32'h00000000,
        RAM[8058] = 32'h00000000,
        RAM[8059] = 32'h00000000,
        RAM[8060] = 32'h00000000,
        RAM[8061] = 32'h00000000,
        RAM[8062] = 32'h00000000,
        RAM[8063] = 32'h00000000,
        RAM[8064] = 32'h00000000,
        RAM[8065] = 32'h00000000,
        RAM[8066] = 32'h00000000,
        RAM[8067] = 32'h00000000,
        RAM[8068] = 32'h00000000,
        RAM[8069] = 32'h00000000,
        RAM[8070] = 32'h00000000,
        RAM[8071] = 32'h00000000,
        RAM[8072] = 32'h00000000,
        RAM[8073] = 32'h00000000,
        RAM[8074] = 32'h00000000,
        RAM[8075] = 32'h00000000,
        RAM[8076] = 32'h00000000,
        RAM[8077] = 32'h00000000,
        RAM[8078] = 32'h00000000,
        RAM[8079] = 32'h00000000,
        RAM[8080] = 32'h00000000,
        RAM[8081] = 32'h00000000,
        RAM[8082] = 32'h00000000,
        RAM[8083] = 32'h00000000,
        RAM[8084] = 32'h00000000,
        RAM[8085] = 32'h00000000,
        RAM[8086] = 32'h00000000,
        RAM[8087] = 32'h00000000,
        RAM[8088] = 32'h00000000,
        RAM[8089] = 32'h00000000,
        RAM[8090] = 32'h00000000,
        RAM[8091] = 32'h00000000,
        RAM[8092] = 32'h00000000,
        RAM[8093] = 32'h00000000,
        RAM[8094] = 32'h00000000,
        RAM[8095] = 32'h00000000,
        RAM[8096] = 32'h00000000,
        RAM[8097] = 32'h00000000,
        RAM[8098] = 32'h00000000,
        RAM[8099] = 32'h00000000,
        RAM[8100] = 32'h00000000,
        RAM[8101] = 32'h00000000,
        RAM[8102] = 32'h00000000,
        RAM[8103] = 32'h00000000,
        RAM[8104] = 32'h00000000,
        RAM[8105] = 32'h00000000,
        RAM[8106] = 32'h00000000,
        RAM[8107] = 32'h00000000,
        RAM[8108] = 32'h00000000,
        RAM[8109] = 32'h00000000,
        RAM[8110] = 32'h00000000,
        RAM[8111] = 32'h00000000,
        RAM[8112] = 32'h00000000,
        RAM[8113] = 32'h00000000,
        RAM[8114] = 32'h00000000,
        RAM[8115] = 32'h00000000,
        RAM[8116] = 32'h00000000,
        RAM[8117] = 32'h00000000,
        RAM[8118] = 32'h00000000,
        RAM[8119] = 32'h00000000,
        RAM[8120] = 32'h00000000,
        RAM[8121] = 32'h00000000,
        RAM[8122] = 32'h00000000,
        RAM[8123] = 32'h00000000,
        RAM[8124] = 32'h00000000,
        RAM[8125] = 32'h00000000,
        RAM[8126] = 32'h00000000,
        RAM[8127] = 32'h00000000,
        RAM[8128] = 32'h00000000,
        RAM[8129] = 32'h00000000,
        RAM[8130] = 32'h00000000,
        RAM[8131] = 32'h00000000,
        RAM[8132] = 32'h00000000,
        RAM[8133] = 32'h00000000,
        RAM[8134] = 32'h00000000,
        RAM[8135] = 32'h00000000,
        RAM[8136] = 32'h00000000,
        RAM[8137] = 32'h00000000,
        RAM[8138] = 32'h00000000,
        RAM[8139] = 32'h00000000,
        RAM[8140] = 32'h00000000,
        RAM[8141] = 32'h00000000,
        RAM[8142] = 32'h00000000,
        RAM[8143] = 32'h00000000,
        RAM[8144] = 32'h00000000,
        RAM[8145] = 32'h00000000,
        RAM[8146] = 32'h00000000,
        RAM[8147] = 32'h00000000,
        RAM[8148] = 32'h00000000,
        RAM[8149] = 32'h00000000,
        RAM[8150] = 32'h00000000,
        RAM[8151] = 32'h00000000,
        RAM[8152] = 32'h00000000,
        RAM[8153] = 32'h00000000,
        RAM[8154] = 32'h00000000,
        RAM[8155] = 32'h00000000,
        RAM[8156] = 32'h00000000,
        RAM[8157] = 32'h00000000,
        RAM[8158] = 32'h00000000,
        RAM[8159] = 32'h00000000,
        RAM[8160] = 32'h00000000,
        RAM[8161] = 32'h00000000,
        RAM[8162] = 32'h00000000,
        RAM[8163] = 32'h00000000,
        RAM[8164] = 32'h00000000,
        RAM[8165] = 32'h00000000,
        RAM[8166] = 32'h00000000,
        RAM[8167] = 32'h00000000,
        RAM[8168] = 32'h00000000,
        RAM[8169] = 32'h00000000,
        RAM[8170] = 32'h00000000,
        RAM[8171] = 32'h00000000,
        RAM[8172] = 32'h00000000,
        RAM[8173] = 32'h00000000,
        RAM[8174] = 32'h00000000,
        RAM[8175] = 32'h00000000,
        RAM[8176] = 32'h00000000,
        RAM[8177] = 32'h00000000,
        RAM[8178] = 32'h00000000,
        RAM[8179] = 32'h00000000,
        RAM[8180] = 32'h00000000,
        RAM[8181] = 32'h00000000,
        RAM[8182] = 32'h00000000,
        RAM[8183] = 32'h00000000,
        RAM[8184] = 32'h00000000,
        RAM[8185] = 32'h00000000,
        RAM[8186] = 32'h00000000,
        RAM[8187] = 32'h00000000,
        RAM[8188] = 32'h00000000,
        RAM[8189] = 32'h00000000,
        RAM[8190] = 32'h00000000,
        RAM[8191] = 32'h00000000,
    end

    always @ (posedge clk)begin
        if(ena == 1)begin
              if(wea[0] == 1)begin
                 douta[7:0] <= dina[7:0];
                 RAM[addra[data_mem_size_in_bits-1:2]][7:0] <= dina[7:0];
              end
              else begin
                 douta[7:0] <= RAM[addra[data_mem_size_in_bits-1:2]][7:0]
              end

              if(wea[1] == 1)begin
                 douta[15:8] <= dina[15:8];
                 RAM[addra[data_mem_size_in_bits-1:2]][15:8] <= dina[15:8]
              end
              else begin
                 douta[15:8] <= RAM[addra[data_mem_size_in_bits-1:2]][15:8];
              end

              if(wea[2] == 1)begin
                 douta[23:16] <= dina[23:16];
                 RAM[addra[data_mem_size_in_bits-1:2]][23:16] <= dina[23:16];
              end
              else begin
                 douta[23:16] <= RAM[addra[data_mem_size_in_bits-1:2]][23:16]; 
              end

              if(wea[3] == 1)begin
                 douta[31:24] <= dina[31:24];
                 RAM[addra[data_mem_size_in_bits-1:2]][31:24] <= dina[31:24];
              end
              else begin
                 douta[31:24] <= RAM[addra[data_mem_size_in_bits-1:2]][31:24];
              end

        end
   end

    always @ (posedge clk)begin
        if(enb == 1)begin
              if(web[0] == 1)begin
                 doutb[7:0] <= dinb[7:0];
                 RAM[addrb[data_mem_size_in_bits-1:2]][7:0] <= dinb[7:0];
              end
              else begin
                 doutb[7:0] <= RAM[addrb[data_mem_size_in_bits-1:2]][7:0]
              end

              if(web[1] == 1)begin
                 doutb[15:8] <= dinb[15:8];
                 RAM[addrb[data_mem_size_in_bits-1:2]][15:8] <= dinb[15:8]
              end
              else begin
                 doutb[15:8] <= RAM[addrb[data_mem_size_in_bits-1:2]][15:8];
              end

              if(web[2] == 1)begin
                 doutb[23:16] <= dinb[23:16];
                 RAM[addrb[data_mem_size_in_bits-1:2]][23:16] <= dinb[23:16];
              end
              else begin
                 doutb[23:16] <= RAM[addrb[data_mem_size_in_bits-1:2]][23:16]; 
              end

              if(web[3] == 1)begin
                 doutb[31:24] <= dinb[31:24];
                 RAM[addrb[data_mem_size_in_bits-1:2]][31:24] <= dinb[31:24];
              end
              else begin
                 doutb[31:24] <= RAM[addrb[data_mem_size_in_bits-1:2]][31:24];
              end

        end
   end
endmodule
